module add
(input wire add,
input wire sub,
input wire div,
input wire mul,
input wire pow,
input wire act_func,
input wire act_func_2_1,

	 input wire[16:0] r1,
	 input wire[16:0] r2,
	 output wire[32:0] output_reg
);
reg[224:0] data;
always @(add, sub, div, mul, pow, act_func, act_func_2_1, r1,r2)
begin
case ({r1, r2})
32'b00000000000000010000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111011;
32'b00000000000000010000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000111111;
32'b00000000000000010000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000111111;
32'b00000000000000010000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000111111;
32'b00000000000000010000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111;
32'b00000000000000010000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000111111;
32'b00000000000000010000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000111111;
32'b00000000000000010000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000111111;
32'b00000000000000010000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000010100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000011000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000000100000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011000010011;
32'b00000000000000100000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000101000101011;
32'b00000000000000100000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000001000101011;
32'b00000000000000100000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000001000101011;
32'b00000000000000100000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000001000101011;
32'b00000000000000100000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000001000101011;
32'b00000000000000100000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000001000101011;
32'b00000000000000100000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000001000101011;
32'b00000000000000100000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000100100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101011;
32'b00000000000000101000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001101011;
32'b00000000000001000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000010011;
32'b00000000000001000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001010001010000000011;
32'b00000000000001000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000010101000000000000000000000000101011;
32'b00000000000001000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000010000000000010000100000000000000000000000000000000000101011;
32'b00000000000001000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000101111;
32'b00000000000001000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011110110000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000101111;
32'b00000000000001000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000101111;
32'b00000000000001000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000101111;
32'b00000000000001000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000001000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000101111;
32'b00000000000001000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000101111;
32'b00000000000001000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111;
32'b00000000000001000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000101111;
32'b00000000000001000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011111000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000101111;
32'b00000000000001000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001101111;
32'b00000000000001001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101111;
32'b00000000000010000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000000000001000010011;
32'b00000000000010000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000010000000010100010000000010000000011;
32'b00000000000010000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000100000000000000000010000100000000000000000000000000001010000000011;
32'b00000000000010000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110000000000000000000000000000000010000000000010000000000000000001000000000000000000000000000000000000000000101011;
32'b00000000000010000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000001000101011;
32'b00000000000010000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011110110010000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000101011;
32'b00000000000010000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000001000000000000101011;
32'b00000000000010000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000010010000000000000000000000000000000000001000000000000000000000000000000000101011;
32'b00000000000010000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000001000101011;
32'b00000000000010000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000000000000000001000000001000000000000000000000000000000000000000000000000000000000100000000000000000101011;
32'b00000000000010000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000001000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000101011;
32'b00000000000010000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000011010110000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000101011;
32'b00000000000010000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000011010111000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000101011;
32'b00000000000010000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100010001010110000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000001101011;
32'b00000000000010000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000100000001010110000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000010000000101011;
32'b00000000000010001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100100000001010110000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000100000000000000101011;
32'b00000000000100000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000000000001000010011;
32'b00000000000100000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000100000000101000100000000100000000000000011;
32'b00000000000100000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000010000000010000000111;
32'b00000000000100000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000001010000000111;
32'b00000000000100000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111111;
32'b00000000000100000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000101111;
32'b00000000000100000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000101111;
32'b00000000000100000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000101111;
32'b00000000000100000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000000100000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000101111;
32'b00000000000100000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000101111;
32'b00000000000100000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011111000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000101111;
32'b00000000000100000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111;
32'b00000000000100000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000101111;
32'b00000000000100000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000101111;
32'b00000000000100001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000101111;
32'b00000000001000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000110100000000000000000000000000001000010011;
32'b00000000001000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000001000000001010001000000000000000100000000000000011;
32'b00000000001000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110110000000000000000000000000000000000000100000000100000000010000000000000000000000000000100000000000000010000000011;
32'b00000000001000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011110110010000000000000001000000000000000000000000000000100000000000000000000000000000000000000000010000000010000000011;
32'b00000000001000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000011010110000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000001011000000011;
32'b00000000001000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000011010110000000000000000000000000000000000010000000010000000000000000000000000000010000000000000000000000000000000101011;
32'b00000000001000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000001000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000101011;
32'b00000000001000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000000000000001001000000000000000000000000000000000000000000000000000000000000000010000000000000000000101011;
32'b00000000001000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000101011;
32'b00000000001000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000100000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101011;
32'b00000000001000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000011010111000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000101011;
32'b00000000001000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000001101011;
32'b00000000001000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010001000101011;
32'b00000000001000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110110000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000100000101011;
32'b00000000001000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000001110110000000000000000000000000000000000000000000000100000000000000000010000000000000000001000000000000000000000101011;
32'b00000000001000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000001000000000001000000000000000000000000000000000000000000000010000000000000000000000000000101011;
32'b00000000010000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000001101000000000000000000000000000000000001000010011;
32'b00000000010000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000010000000010100010000000000000001000000000000000000000011;
32'b00000000010000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011110110000000000000000000000010000000000000000000000000100000000000000000000000000001001000000000000100000000000000011;
32'b00000000010000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000000000000000000000000001000000000010000000000000000000000000000000100000001000000010000000011;
32'b00000000010000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000010000000010000000111;
32'b00000000010000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001010000000111;
32'b00000000010000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000101111;
32'b00000000010000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000101111;
32'b00000000010000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011011110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
32'b00000000010000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011011111000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111;
32'b00000000010000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001101111;
32'b00000000010000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000101111;
32'b00000000010000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000101111;
32'b00000000010000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000101111;
32'b00000000010000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000101111;
32'b00000000010000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000101111;
32'b00000000100000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000011010000000000000000000000000000000000000000001000010011;
32'b00000000100000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000100000000101000100000000000000000000001000000000000000000000011;
32'b00000000100000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011110110000000001000000000000000000000000000000001000000000000000000000000000010000000000000000000000100000001000000011;
32'b00000000100000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000000000000000000010000000000000000000000001000000000001000001000000000000000000000010000000011;
32'b00000000100000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000000000000000000010000100000000000000000000000000000000000000000000000000000000100000000000000011000000011;
32'b00000000100000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000000000000000001000000000000000000000000000000000000001000000000000000000000000010000010000000010000000011;
32'b00000000100000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010011010110000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000001011000000011;
32'b00000000100000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000011010110000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000101011;
32'b00000000100000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011011111000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000101011;
32'b00000000100000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001101011;
32'b00000000100000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000001110110000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010001000101011;
32'b00000000100000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110110000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000100000000000000101011;
32'b00000000100000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101000001010110000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000001000101011;
32'b00000000100000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101000001010110000000000000000000000000000001000000000000000000000000000001000000000000000010000000000000000000000000000101011;
32'b00000000100000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100010001010110000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000001000101011;
32'b00000000100000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000100000001010110000000000000000000000000000000000000000000010000000000000001001000000000000000000000000000000000000000000101011;
32'b00000001000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000110100000000000000000000000000000000000000000000000001000010011;
32'b00000001000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000001000000001010001000000000000000000000010000000000000000000000000000011;
32'b00000001000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000100000000000010111;
32'b00000001000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011011110000000000000000000000000000100000000000000000000001000000000000000000010000000000000000000000100000000000000111;
32'b00000001000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000010000010111;
32'b00000001000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011110000000000000010000000000000000000000000000000000001000000000000000000000000000000000100000000000000010000000111;
32'b00000001000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011011110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000010111;
32'b00000001000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011011111000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001010000000111;
32'b00000001000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111;
32'b00000001000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000101111;
32'b00000001000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000111111;
32'b00000001000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000101111;
32'b00000001000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111;
32'b00000001000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000101111;
32'b00000001000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000111111;
32'b00000001000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000101111;
32'b00000010000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000001101000000000000000000000000000000000000000000000000000000001000010011;
32'b00000010000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000010000000010100010000000000000000000000000000010000000000000000000000000000011;
32'b00000010000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000000000000100000000000000000000000000001000000000000000000000000000001000001000000001000000011;
32'b00000010000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000000000000000001000000001000000000000000100000000000000000100000000000000000000000000000100000000000000011;
32'b00000010000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000000000010000000000000000000000000000000000000000000000000000000010000000100000000000000000000011000000011;
32'b00000010000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000011010110000000100000000100000000000000000000000000000100000000000000000000000000000001000000000000000000000010000000011;
32'b00000010000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000011010111000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000011000000011;
32'b00000010000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000001010110010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000010001000011;
32'b00000010000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000011011000000011;
32'b00000010000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000100000101011;
32'b00000010000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001010110000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000001000101011;
32'b00000010000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100010001010110000000000000000000000000000000000000000000000100000000000000000000000000000010000000010000000000000000000101011;
32'b00000010000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100100000001010110000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000001000101011;
32'b00000010000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100100000001010110000000000000000000000000000000000000000000000100000000000000001000000001000000000000000000000000000000000101011;
32'b00000010000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000001010110000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000101011;
32'b00000010000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000001110110000000000000000000000000000000000000000000000100100000000100000000000000000000000000000000000000000000000101011;
32'b00000100000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000011010000000000000000000000000000000000000000000000000000000000000001000010011;
32'b00000100000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000100000000101000100000000000000000000000000000100000000000000000000000000000000000011;
32'b00000100000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000000000000000001000000000000000000000000000010000000000000000000000000000101000001000000000000000000000011;
32'b00000100000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010110000000001000010000000000000000000000000000000000000010001000000000000000000000000000000000000100000000000000011;
32'b00000100000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010011010110000000100000000000000000000000000000000000000000001000000000000100000000000000000000000000000100000000000000111;
32'b00000100000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000011010111000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000010000000111;
32'b00000100000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000010001000111;
32'b00000100000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000010010000000111;
32'b00000100000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010000010111;
32'b00000100000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000001010000000111;
32'b00000100000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000101111;
32'b00000100000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000101111;
32'b00000100000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000101111;
32'b00000100000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000101111;
32'b00000100000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000101111;
32'b00000100000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000101111;
32'b00001000000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000001000010011;
32'b00001000000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000001000000001010001000000000000000000000000000000000000100000000000000000000000000000000000011;
32'b00001000000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000011010110000000000000010000000000000000000000000000100100000000000000000010000000000000000000001000000000000000000000011;
32'b00001000000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000011010110000000100000000000000000000000000000000000000000010000000000000000000000000000000000000100000100000100000000011;
32'b00001000000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000011010111000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000100000001000000011;
32'b00001000000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000000000000010000000000000000000000000100000100000000000000000000000000000000000010001000011;
32'b00001000000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000001110110000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000001000010010000000011;
32'b00001000000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000100000000000000000000000000000000000000000000000000000000000001000000000100100000000010000000011;
32'b00001000000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101000001010110000000000000000000000000000000000000000000000000001000000000000000000000000000000001100000000000000011000000011;
32'b00001000000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100100000001010110000000000000000000000000000000010000000000000000000000000000000000000000000010000000010000010000000010000000011;
32'b00001000000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100010001010110000000001000000000000000000000000000000000000100000000000000000000000100000000000000000000000000001010000000011;
32'b00001000000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000000000000000000000000010000000000000000001000000000000000000000000100000000000000000101011;
32'b00001000000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110110000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000001000101011;
32'b00001000000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000001110110010000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000101011;
32'b00001000000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000100001000100000000000000000000000000000000000000000000000000000000000101011;
32'b00001000000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100100000001010110000000000000000000000000000000000010000000000000000000000000000000000001000000000000000100000000000000000101011;
32'b00010000000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000001000010011;
32'b00010000000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000010000000010100010000000000000000000000000000000000001000000000000000000000000000000000000000000011;
32'b00010000000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011010110000000100000000000000000000000000001000000000000001000000000000000000000000000010000000000000000000000000000111;
32'b00010000000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011011111000000000000000000000000000000000000000000100000000000000000000000000000000000100000001000000000000000000000111;
32'b00010000000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000001010111;
32'b00010000000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000100010000000000111;
32'b00010000000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000100000000010000000111;
32'b00010000000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000000000000000000000000010000000100001000000000000000010000000111;
32'b00010000000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000010000010111;
32'b00010000000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000010000000000000000000000000000000000000000000000100000000000000100000000000000010000000111;
32'b00010000000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000010000000010000000111;
32'b00010000000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000001010000000111;
32'b00010000000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111111;
32'b00010000000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000101111;
32'b00010000000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000101111;
32'b00010000000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000101111;
32'b00100000000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011;
32'b00100000000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000100000000101000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000011;
32'b00100000000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000011010111000000000000000000000000000010000000100000000100000000000000000000000000000000010000000000000000000000000000011;
32'b00100000000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100010001010110000000000000000000000000000000000001000000000000000000000100000000000000010000000000001000000000000000001000011;
32'b00100000000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000100010001000000011;
32'b00100000000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110110000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000100100000100000000011;
32'b00100000000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000001110110000000001000000000000000000000000000000000000100000000001000000000000000000000000001000000000000000010000000011;
32'b00100000000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101000001010110000000000000000000000000000001000000000000000000000000000000000100000000010010000000000000000000000010000000011;
32'b00100000000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100100000001010110000000000000000000000000000000000000000000000000001000000000000000000110000000000000000000000000000011000000011;
32'b00100000000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100100000001010110000000000000000001000000000000000000000000000000000000000000001000000001000001000000000000000000000010000000011;
32'b00100000000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000000000000000000000000000100000000010000000000000000000000000000100000001000000010000000011;
32'b00100000000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000001110110010000000000000000000000000000000000000000000000100000000000000000000000010000000000000000010000000010000000011;
32'b00100000000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101000001010110000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000001011000000011;
32'b00100000000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000100000001010110000000000000000001000000000000000010000000010000000000000000000000000000000000000000000000000000000000000101011;
32'b00100000000000000100000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000000000100000000000000000100000000000000000010000000000000000000000000000000000000000101011;
32'b00100000000000001000000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000001000000000000000000000000000000010000000000000000000000000000000010000000000000000000101011;
32'b01000000000000000000000000000001: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011;
32'b01000000000000000000000000000010: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011;
32'b01000000000000000000000000000100: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000001000011;
32'b01000000000000000000000000001000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000100000001010110000000000000000000000000000010000000100000000000000010000000000000000000000000000000001000000000010000000000011;
32'b01000000000000000000000000010000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001010110000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000100100000000000000111;
32'b01000000000000000000000000100000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000001110110000000000000000000000000000000000000000000100000000000000000000010000000000000000001000000000100000000000000111;
32'b01000000000000000000000001000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000000000000000010000000000000000000000000010100000000000000100000000000000111;
32'b01000000000000000000000010000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000001000000010000000111;
32'b01000000000000000000000100000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000010000010111;
32'b01000000000000000000001000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000001000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000010000000111;
32'b01000000000000000000010000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111110000000000000000000000010000000000000000000000000100000000000000000000000000001000000000000000000000010000000111;
32'b01000000000000000000100000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001011110000000000000000000000000000000000000100001000000000000000000000000000000000000000000100000000000000010000000111;
32'b01000000000000000001000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001011110000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000010000000010000000111;
32'b01000000000000000010000000000000: data <= 224'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011110000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000001010000000111;
module add
(input wire add,
input wire sub,
input wire div,
input wire mul,
input wire pow,
input wire act_func,
input wire act_func_2_1,

	 input wire[16:0] r1,
	 input wire[16:0] r2,
	 output wire[32:0] output_reg
);
assign output_reg = {r1[3]&r2[5]&pow|r1[3]&r2[11]&pow|r1[3]&r2[12]&pow|r1[3]&r2[14]&pow|r1[4]&r2[12]&div|r1[4]&r2[13]&div|r1[4]&r2[14]&div|r1[4]&r2[15]&div|r1[5]&r2[3]&pow|r1[5]&r2[4]&pow|r1[5]&r2[5]&pow|r1[5]&r2[10]&div|r1[5]&r2[10]&pow|r1[5]&r2[11]&div|r1[5]&r2[12]&div|r1[6]&r2[8]&div|r1[6]&r2[9]&div|r1[6]&r2[10]&div|r1[7]&r2[2]&pow|r1[7]&r2[7]&div|r1[7]&r2[7]&pow|r1[7]&r2[8]&div|r1[7]&r2[9]&div|r1[7]&r2[10]&pow|r1[7]&r2[15]&pow|r1[8]&r2[6]&div|r1[8]&r2[7]&div|r1[8]&r2[14]&div|r1[8]&r2[15]&div|r1[9]&r2[6]&div|r1[9]&r2[6]&pow|r1[9]&r2[7]&div|r1[9]&r2[7]&pow|r1[9]&r2[13]&div|r1[9]&r2[14]&div|r1[9]&r2[14]&pow|r1[9]&r2[15]&pow|r1[10]&r2[5]&div|r1[10]&r2[6]&div|r1[10]&r2[12]&div|r1[11]&r2[2]&pow|r1[11]&r2[3]&pow|r1[11]&r2[4]&pow|r1[11]&r2[5]&div|r1[11]&r2[11]&div|r1[11]&r2[13]&pow|r1[12]&r2[4]&div|r1[12]&r2[5]&div|r1[12]&r2[10]&div|r1[12]&r2[15]&div|r1[13]&r2[4]&div|r1[13]&r2[6]&pow|r1[13]&r2[9]&div|r1[13]&r2[11]&pow|r1[13]&r2[12]&pow|r1[13]&r2[13]&pow|r1[13]&r2[14]&div|r1[14]&r2[3]&pow|r1[14]&r2[4]&div|r1[14]&r2[8]&div|r1[14]&r2[9]&div|r1[14]&r2[13]&div|r1[15]&r2[4]&div|r1[15]&r2[8]&div|r1[15]&r2[12]&div,
r1[2]&r2[5]&pow|r1[3]&r2[8]&pow|r1[3]&r2[9]&pow|r1[3]&r2[10]&pow|r1[3]&r2[11]&div|r1[3]&r2[12]&div|r1[3]&r2[13]&div|r1[3]&r2[14]&div|r1[3]&r2[15]&div|r1[3]&r2[15]&pow|r1[4]&r2[8]&div|r1[4]&r2[9]&div|r1[4]&r2[10]&div|r1[4]&r2[11]&div|r1[5]&r2[7]&div|r1[5]&r2[7]&pow|r1[5]&r2[8]&div|r1[5]&r2[8]&pow|r1[5]&r2[9]&div|r1[5]&r2[9]&pow|r1[5]&r2[14]&pow|r1[6]&r2[2]&pow|r1[6]&r2[5]&pow|r1[6]&r2[6]&div|r1[6]&r2[7]&div|r1[7]&r2[4]&pow|r1[7]&r2[5]&div|r1[7]&r2[5]&pow|r1[7]&r2[6]&div|r1[7]&r2[12]&pow|r1[7]&r2[13]&pow|r1[7]&r2[14]&div|r1[7]&r2[15]&div|r1[8]&r2[4]&div|r1[8]&r2[5]&div|r1[8]&r2[12]&div|r1[8]&r2[13]&div|r1[9]&r2[4]&div|r1[9]&r2[4]&pow|r1[9]&r2[5]&div|r1[9]&r2[5]&pow|r1[9]&r2[11]&div|r1[9]&r2[12]&div|r1[9]&r2[12]&pow|r1[9]&r2[13]&pow|r1[10]&r2[2]&pow|r1[10]&r2[3]&pow|r1[10]&r2[4]&div|r1[10]&r2[5]&pow|r1[10]&r2[10]&div|r1[10]&r2[11]&div|r1[11]&r2[3]&div|r1[11]&r2[4]&div|r1[11]&r2[6]&pow|r1[11]&r2[8]&pow|r1[11]&r2[9]&div|r1[11]&r2[9]&pow|r1[11]&r2[10]&div|r1[11]&r2[15]&div|r1[11]&r2[15]&pow|r1[12]&r2[3]&div|r1[12]&r2[8]&div|r1[12]&r2[9]&div|r1[12]&r2[14]&div|r1[13]&r2[2]&pow|r1[13]&r2[3]&div|r1[13]&r2[7]&pow|r1[13]&r2[8]&div|r1[13]&r2[8]&pow|r1[13]&r2[9]&pow|r1[13]&r2[13]&div|r1[14]&r2[3]&div|r1[14]&r2[5]&pow|r1[14]&r2[7]&div|r1[14]&r2[12]&div|r1[15]&r2[2]&pow|r1[15]&r2[3]&div|r1[15]&r2[3]&pow|r1[15]&r2[6]&pow|r1[15]&r2[7]&div|r1[15]&r2[7]&pow|r1[15]&r2[10]&pow|r1[15]&r2[11]&div|r1[15]&r2[11]&pow|r1[15]&r2[14]&pow|r1[15]&r2[15]&div,
r1[1]&r2[15]&add|r1[2]&r2[4]&pow|r1[2]&r2[8]&div|r1[2]&r2[9]&div|r1[2]&r2[10]&div|r1[2]&r2[11]&div|r1[2]&r2[12]&div|r1[2]&r2[13]&div|r1[2]&r2[14]&add|r1[2]&r2[14]&div|r1[2]&r2[15]&add|r1[2]&r2[15]&div|r1[3]&r2[3]&pow|r1[3]&r2[4]&pow|r1[3]&r2[6]&div|r1[3]&r2[6]&pow|r1[3]&r2[7]&div|r1[3]&r2[8]&div|r1[3]&r2[9]&div|r1[3]&r2[10]&div|r1[3]&r2[13]&add|r1[3]&r2[13]&pow|r1[3]&r2[14]&add|r1[3]&r2[15]&add|r1[4]&r2[2]&pow|r1[4]&r2[4]&div|r1[4]&r2[5]&div|r1[4]&r2[6]&div|r1[4]&r2[7]&div|r1[4]&r2[12]&add|r1[4]&r2[13]&add|r1[4]&r2[14]&add|r1[4]&r2[15]&add|r1[5]&r2[2]&pow|r1[5]&r2[4]&div|r1[5]&r2[5]&div|r1[5]&r2[6]&div|r1[5]&r2[11]&add|r1[5]&r2[11]&pow|r1[5]&r2[12]&add|r1[5]&r2[12]&pow|r1[5]&r2[13]&add|r1[5]&r2[13]&pow|r1[5]&r2[14]&add|r1[5]&r2[15]&add|r1[6]&r2[3]&div|r1[6]&r2[3]&pow|r1[6]&r2[4]&div|r1[6]&r2[4]&pow|r1[6]&r2[5]&div|r1[6]&r2[10]&add|r1[6]&r2[11]&add|r1[6]&r2[12]&add|r1[6]&r2[13]&add|r1[6]&r2[14]&add|r1[6]&r2[14]&div|r1[6]&r2[15]&add|r1[6]&r2[15]&div|r1[7]&r2[3]&div|r1[7]&r2[3]&pow|r1[7]&r2[4]&div|r1[7]&r2[6]&pow|r1[7]&r2[9]&add|r1[7]&r2[10]&add|r1[7]&r2[11]&add|r1[7]&r2[11]&pow|r1[7]&r2[12]&add|r1[7]&r2[12]&div|r1[7]&r2[13]&add|r1[7]&r2[13]&div|r1[7]&r2[14]&add|r1[7]&r2[14]&pow|r1[7]&r2[15]&add|r1[8]&r2[2]&div|r1[8]&r2[3]&div|r1[8]&r2[8]&add|r1[8]&r2[9]&add|r1[8]&r2[10]&add|r1[8]&r2[10]&div|r1[8]&r2[11]&add|r1[8]&r2[11]&div|r1[8]&r2[12]&add|r1[8]&r2[13]&add|r1[8]&r2[14]&add|r1[8]&r2[15]&add|r1[9]&r2[2]&div|r1[9]&r2[2]&pow|r1[9]&r2[3]&div|r1[9]&r2[3]&pow|r1[9]&r2[7]&add|r1[9]&r2[8]&add|r1[9]&r2[9]&add|r1[9]&r2[9]&div|r1[9]&r2[10]&add|r1[9]&r2[10]&div|r1[9]&r2[10]&pow|r1[9]&r2[11]&add|r1[9]&r2[11]&pow|r1[9]&r2[12]&add|r1[9]&r2[13]&add|r1[9]&r2[14]&add|r1[9]&r2[15]&add|r1[10]&r2[2]&div|r1[10]&r2[3]&div|r1[10]&r2[4]&pow|r1[10]&r2[6]&add|r1[10]&r2[7]&add|r1[10]&r2[8]&add|r1[10]&r2[8]&div|r1[10]&r2[9]&add|r1[10]&r2[9]&div|r1[10]&r2[10]&add|r1[10]&r2[11]&add|r1[10]&r2[12]&add|r1[10]&r2[13]&add|r1[10]&r2[14]&add|r1[10]&r2[15]&add|r1[10]&r2[15]&div|r1[11]&r2[2]&div|r1[11]&r2[5]&add|r1[11]&r2[5]&pow|r1[11]&r2[6]&add|r1[11]&r2[7]&add|r1[11]&r2[8]&add|r1[11]&r2[8]&div|r1[11]&r2[9]&add|r1[11]&r2[10]&add|r1[11]&r2[10]&pow|r1[11]&r2[11]&add|r1[11]&r2[11]&pow|r1[11]&r2[12]&add|r1[11]&r2[12]&pow|r1[11]&r2[13]&add|r1[11]&r2[14]&add|r1[11]&r2[14]&div|r1[11]&r2[15]&add|r1[12]&r2[2]&div|r1[12]&r2[2]&pow|r1[12]&r2[4]&add|r1[12]&r2[5]&add|r1[12]&r2[6]&add|r1[12]&r2[7]&add|r1[12]&r2[7]&div|r1[12]&r2[8]&add|r1[12]&r2[9]&add|r1[12]&r2[10]&add|r1[12]&r2[11]&add|r1[12]&r2[12]&add|r1[12]&r2[12]&div|r1[12]&r2[13]&add|r1[12]&r2[13]&div|r1[12]&r2[14]&add|r1[12]&r2[15]&add|r1[13]&r2[2]&div|r1[13]&r2[3]&add|r1[13]&r2[3]&pow|r1[13]&r2[4]&add|r1[13]&r2[4]&pow|r1[13]&r2[5]&add|r1[13]&r2[5]&pow|r1[13]&r2[6]&add|r1[13]&r2[7]&add|r1[13]&r2[7]&div|r1[13]&r2[8]&add|r1[13]&r2[9]&add|r1[13]&r2[10]&add|r1[13]&r2[11]&add|r1[13]&r2[12]&add|r1[13]&r2[12]&div|r1[13]&r2[13]&add|r1[13]&r2[14]&add|r1[13]&r2[14]&pow|r1[13]&r2[15]&add|r1[14]&r2[2]&add|r1[14]&r2[2]&div|r1[14]&r2[3]&add|r1[14]&r2[4]&add|r1[14]&r2[4]&pow|r1[14]&r2[5]&add|r1[14]&r2[6]&add|r1[14]&r2[6]&div|r1[14]&r2[7]&add|r1[14]&r2[8]&add|r1[14]&r2[9]&add|r1[14]&r2[10]&add|r1[14]&r2[11]&add|r1[14]&r2[11]&div|r1[14]&r2[12]&add|r1[14]&r2[13]&add|r1[14]&r2[14]&add|r1[14]&r2[15]&add|r1[14]&r2[15]&div|r1[15]&r2[1]&add|r1[15]&r2[2]&add|r1[15]&r2[2]&div|r1[15]&r2[3]&add|r1[15]&r2[4]&add|r1[15]&r2[5]&add|r1[15]&r2[6]&add|r1[15]&r2[6]&div|r1[15]&r2[7]&add|r1[15]&r2[8]&add|r1[15]&r2[9]&add|r1[15]&r2[10]&add|r1[15]&r2[10]&div|r1[15]&r2[11]&add|r1[15]&r2[12]&add|r1[15]&r2[13]&add|r1[15]&r2[14]&add|r1[15]&r2[14]&div|r1[15]&r2[15]&add,
r1[0]&r2[0]&add|r1[0]&r2[0]&sub|r1[0]&r2[0]&div|r1[0]&r2[0]&mul|r1[0]&r2[0]&pow|r1[0]&r2[0]&act_func|r1[0]&r2[0]&act_func_2_1|r1[0]&r2[1]&add|r1[0]&r2[1]&sub|r1[0]&r2[1]&div|r1[0]&r2[1]&mul|r1[0]&r2[1]&pow|r1[0]&r2[1]&act_func|r1[0]&r2[1]&act_func_2_1|r1[0]&r2[2]&add|r1[0]&r2[2]&sub|r1[0]&r2[2]&div|r1[0]&r2[2]&mul|r1[0]&r2[2]&pow|r1[0]&r2[2]&act_func|r1[0]&r2[2]&act_func_2_1|r1[0]&r2[3]&add|r1[0]&r2[3]&sub|r1[0]&r2[3]&div|r1[0]&r2[3]&mul|r1[0]&r2[3]&pow|r1[0]&r2[3]&act_func|r1[0]&r2[3]&act_func_2_1|r1[0]&r2[4]&add|r1[0]&r2[4]&sub|r1[0]&r2[4]&div|r1[0]&r2[4]&mul|r1[0]&r2[4]&pow|r1[0]&r2[4]&act_func|r1[0]&r2[4]&act_func_2_1|r1[0]&r2[5]&add|r1[0]&r2[5]&sub|r1[0]&r2[5]&div|r1[0]&r2[5]&mul|r1[0]&r2[5]&pow|r1[0]&r2[5]&act_func|r1[0]&r2[5]&act_func_2_1|r1[0]&r2[6]&add|r1[0]&r2[6]&sub|r1[0]&r2[6]&div|r1[0]&r2[6]&mul|r1[0]&r2[6]&pow|r1[0]&r2[6]&act_func|r1[0]&r2[6]&act_func_2_1|r1[0]&r2[7]&add|r1[0]&r2[7]&sub|r1[0]&r2[7]&div|r1[0]&r2[7]&mul|r1[0]&r2[7]&pow|r1[0]&r2[7]&act_func|r1[0]&r2[7]&act_func_2_1|r1[0]&r2[8]&add|r1[0]&r2[8]&sub|r1[0]&r2[8]&div|r1[0]&r2[8]&mul|r1[0]&r2[8]&pow|r1[0]&r2[8]&act_func|r1[0]&r2[8]&act_func_2_1|r1[0]&r2[9]&add|r1[0]&r2[9]&sub|r1[0]&r2[9]&div|r1[0]&r2[9]&mul|r1[0]&r2[9]&pow|r1[0]&r2[9]&act_func|r1[0]&r2[9]&act_func_2_1|r1[0]&r2[10]&add|r1[0]&r2[10]&sub|r1[0]&r2[10]&div|r1[0]&r2[10]&mul|r1[0]&r2[10]&pow|r1[0]&r2[10]&act_func|r1[0]&r2[10]&act_func_2_1|r1[0]&r2[11]&add|r1[0]&r2[11]&sub|r1[0]&r2[11]&div|r1[0]&r2[11]&mul|r1[0]&r2[11]&pow|r1[0]&r2[11]&act_func|r1[0]&r2[11]&act_func_2_1|r1[0]&r2[12]&add|r1[0]&r2[12]&sub|r1[0]&r2[12]&div|r1[0]&r2[12]&mul|r1[0]&r2[12]&pow|r1[0]&r2[12]&act_func|r1[0]&r2[12]&act_func_2_1|r1[0]&r2[13]&add|r1[0]&r2[13]&sub|r1[0]&r2[13]&div|r1[0]&r2[13]&mul|r1[0]&r2[13]&pow|r1[0]&r2[13]&act_func|r1[0]&r2[13]&act_func_2_1|r1[0]&r2[14]&add|r1[0]&r2[14]&sub|r1[0]&r2[14]&div|r1[0]&r2[14]&mul|r1[0]&r2[14]&pow|r1[0]&r2[14]&act_func|r1[0]&r2[14]&act_func_2_1|r1[0]&r2[15]&add|r1[0]&r2[15]&sub|r1[0]&r2[15]&div|r1[0]&r2[15]&mul|r1[0]&r2[15]&pow|r1[0]&r2[15]&act_func|r1[0]&r2[15]&act_func_2_1|r1[1]&r2[0]&add|r1[1]&r2[0]&sub|r1[1]&r2[0]&div|r1[1]&r2[0]&mul|r1[1]&r2[0]&pow|r1[1]&r2[0]&act_func|r1[1]&r2[0]&act_func_2_1|r1[1]&r2[1]&add|r1[1]&r2[1]&sub|r1[1]&r2[1]&div|r1[1]&r2[1]&mul|r1[1]&r2[1]&pow|r1[1]&r2[1]&act_func|r1[1]&r2[1]&act_func_2_1|r1[1]&r2[2]&add|r1[1]&r2[2]&sub|r1[1]&r2[2]&div|r1[1]&r2[2]&mul|r1[1]&r2[2]&pow|r1[1]&r2[2]&act_func|r1[1]&r2[2]&act_func_2_1|r1[1]&r2[3]&add|r1[1]&r2[3]&sub|r1[1]&r2[3]&div|r1[1]&r2[3]&mul|r1[1]&r2[3]&pow|r1[1]&r2[3]&act_func|r1[1]&r2[3]&act_func_2_1|r1[1]&r2[4]&add|r1[1]&r2[4]&sub|r1[1]&r2[4]&div|r1[1]&r2[4]&mul|r1[1]&r2[4]&pow|r1[1]&r2[4]&act_func|r1[1]&r2[4]&act_func_2_1|r1[1]&r2[5]&add|r1[1]&r2[5]&sub|r1[1]&r2[5]&div|r1[1]&r2[5]&mul|r1[1]&r2[5]&pow|r1[1]&r2[5]&act_func|r1[1]&r2[5]&act_func_2_1|r1[1]&r2[6]&add|r1[1]&r2[6]&sub|r1[1]&r2[6]&div|r1[1]&r2[6]&mul|r1[1]&r2[6]&pow|r1[1]&r2[6]&act_func|r1[1]&r2[6]&act_func_2_1|r1[1]&r2[7]&add|r1[1]&r2[7]&sub|r1[1]&r2[7]&div|r1[1]&r2[7]&mul|r1[1]&r2[7]&pow|r1[1]&r2[7]&act_func|r1[1]&r2[7]&act_func_2_1|r1[1]&r2[8]&add|r1[1]&r2[8]&sub|r1[1]&r2[8]&div|r1[1]&r2[8]&mul|r1[1]&r2[8]&pow|r1[1]&r2[8]&act_func|r1[1]&r2[8]&act_func_2_1|r1[1]&r2[9]&add|r1[1]&r2[9]&sub|r1[1]&r2[9]&div|r1[1]&r2[9]&mul|r1[1]&r2[9]&pow|r1[1]&r2[9]&act_func|r1[1]&r2[9]&act_func_2_1|r1[1]&r2[10]&add|r1[1]&r2[10]&sub|r1[1]&r2[10]&div|r1[1]&r2[10]&mul|r1[1]&r2[10]&pow|r1[1]&r2[10]&act_func|r1[1]&r2[10]&act_func_2_1|r1[1]&r2[11]&add|r1[1]&r2[11]&sub|r1[1]&r2[11]&div|r1[1]&r2[11]&mul|r1[1]&r2[11]&pow|r1[1]&r2[11]&act_func|r1[1]&r2[11]&act_func_2_1|r1[1]&r2[12]&add|r1[1]&r2[12]&sub|r1[1]&r2[12]&div|r1[1]&r2[12]&mul|r1[1]&r2[12]&pow|r1[1]&r2[12]&act_func|r1[1]&r2[12]&act_func_2_1|r1[1]&r2[13]&add|r1[1]&r2[13]&sub|r1[1]&r2[13]&div|r1[1]&r2[13]&mul|r1[1]&r2[13]&pow|r1[1]&r2[13]&act_func|r1[1]&r2[13]&act_func_2_1|r1[1]&r2[14]&add|r1[1]&r2[14]&sub|r1[1]&r2[14]&div|r1[1]&r2[14]&mul|r1[1]&r2[14]&pow|r1[1]&r2[14]&act_func|r1[1]&r2[14]&act_func_2_1|r1[1]&r2[15]&sub|r1[1]&r2[15]&div|r1[1]&r2[15]&mul|r1[1]&r2[15]&pow|r1[1]&r2[15]&act_func|r1[1]&r2[15]&act_func_2_1|r1[2]&r2[0]&add|r1[2]&r2[0]&sub|r1[2]&r2[0]&div|r1[2]&r2[0]&mul|r1[2]&r2[0]&pow|r1[2]&r2[0]&act_func|r1[2]&r2[0]&act_func_2_1|r1[2]&r2[1]&add|r1[2]&r2[1]&sub|r1[2]&r2[1]&div|r1[2]&r2[1]&mul|r1[2]&r2[1]&pow|r1[2]&r2[1]&act_func|r1[2]&r2[1]&act_func_2_1|r1[2]&r2[2]&add|r1[2]&r2[2]&sub|r1[2]&r2[2]&div|r1[2]&r2[2]&mul|r1[2]&r2[2]&pow|r1[2]&r2[2]&act_func|r1[2]&r2[2]&act_func_2_1|r1[2]&r2[3]&add|r1[2]&r2[3]&sub|r1[2]&r2[3]&div|r1[2]&r2[3]&mul|r1[2]&r2[3]&pow|r1[2]&r2[3]&act_func|r1[2]&r2[3]&act_func_2_1|r1[2]&r2[4]&add|r1[2]&r2[4]&sub|r1[2]&r2[4]&div|r1[2]&r2[4]&mul|r1[2]&r2[4]&act_func|r1[2]&r2[4]&act_func_2_1|r1[2]&r2[5]&add|r1[2]&r2[5]&sub|r1[2]&r2[5]&div|r1[2]&r2[5]&mul|r1[2]&r2[5]&act_func|r1[2]&r2[5]&act_func_2_1|r1[2]&r2[6]&add|r1[2]&r2[6]&sub|r1[2]&r2[6]&div|r1[2]&r2[6]&mul|r1[2]&r2[6]&pow|r1[2]&r2[6]&act_func|r1[2]&r2[6]&act_func_2_1|r1[2]&r2[7]&add|r1[2]&r2[7]&sub|r1[2]&r2[7]&div|r1[2]&r2[7]&mul|r1[2]&r2[7]&pow|r1[2]&r2[7]&act_func|r1[2]&r2[7]&act_func_2_1|r1[2]&r2[8]&add|r1[2]&r2[8]&sub|r1[2]&r2[8]&mul|r1[2]&r2[8]&pow|r1[2]&r2[8]&act_func|r1[2]&r2[8]&act_func_2_1|r1[2]&r2[9]&add|r1[2]&r2[9]&sub|r1[2]&r2[9]&mul|r1[2]&r2[9]&pow|r1[2]&r2[9]&act_func|r1[2]&r2[9]&act_func_2_1|r1[2]&r2[10]&add|r1[2]&r2[10]&sub|r1[2]&r2[10]&mul|r1[2]&r2[10]&pow|r1[2]&r2[10]&act_func|r1[2]&r2[10]&act_func_2_1|r1[2]&r2[11]&add|r1[2]&r2[11]&sub|r1[2]&r2[11]&mul|r1[2]&r2[11]&pow|r1[2]&r2[11]&act_func|r1[2]&r2[11]&act_func_2_1|r1[2]&r2[12]&add|r1[2]&r2[12]&sub|r1[2]&r2[12]&mul|r1[2]&r2[12]&pow|r1[2]&r2[12]&act_func|r1[2]&r2[12]&act_func_2_1|r1[2]&r2[13]&add|r1[2]&r2[13]&sub|r1[2]&r2[13]&mul|r1[2]&r2[13]&pow|r1[2]&r2[13]&act_func|r1[2]&r2[13]&act_func_2_1|r1[2]&r2[14]&sub|r1[2]&r2[14]&mul|r1[2]&r2[14]&pow|r1[2]&r2[14]&act_func|r1[2]&r2[14]&act_func_2_1|r1[2]&r2[15]&sub|r1[2]&r2[15]&mul|r1[2]&r2[15]&pow|r1[2]&r2[15]&act_func|r1[2]&r2[15]&act_func_2_1|r1[3]&r2[0]&add|r1[3]&r2[0]&sub|r1[3]&r2[0]&div|r1[3]&r2[0]&mul|r1[3]&r2[0]&pow|r1[3]&r2[0]&act_func|r1[3]&r2[0]&act_func_2_1|r1[3]&r2[1]&add|r1[3]&r2[1]&sub|r1[3]&r2[1]&div|r1[3]&r2[1]&mul|r1[3]&r2[1]&pow|r1[3]&r2[1]&act_func|r1[3]&r2[1]&act_func_2_1|r1[3]&r2[2]&add|r1[3]&r2[2]&sub|r1[3]&r2[2]&div|r1[3]&r2[2]&mul|r1[3]&r2[2]&pow|r1[3]&r2[2]&act_func|r1[3]&r2[2]&act_func_2_1|r1[3]&r2[3]&add|r1[3]&r2[3]&sub|r1[3]&r2[3]&div|r1[3]&r2[3]&mul|r1[3]&r2[3]&act_func|r1[3]&r2[3]&act_func_2_1|r1[3]&r2[4]&add|r1[3]&r2[4]&sub|r1[3]&r2[4]&div|r1[3]&r2[4]&mul|r1[3]&r2[4]&act_func|r1[3]&r2[4]&act_func_2_1|r1[3]&r2[5]&add|r1[3]&r2[5]&sub|r1[3]&r2[5]&div|r1[3]&r2[5]&mul|r1[3]&r2[5]&act_func|r1[3]&r2[5]&act_func_2_1|r1[3]&r2[6]&add|r1[3]&r2[6]&sub|r1[3]&r2[6]&mul|r1[3]&r2[6]&act_func|r1[3]&r2[6]&act_func_2_1|r1[3]&r2[7]&add|r1[3]&r2[7]&sub|r1[3]&r2[7]&mul|r1[3]&r2[7]&pow|r1[3]&r2[7]&act_func|r1[3]&r2[7]&act_func_2_1|r1[3]&r2[8]&add|r1[3]&r2[8]&sub|r1[3]&r2[8]&mul|r1[3]&r2[8]&act_func|r1[3]&r2[8]&act_func_2_1|r1[3]&r2[9]&add|r1[3]&r2[9]&sub|r1[3]&r2[9]&mul|r1[3]&r2[9]&act_func|r1[3]&r2[9]&act_func_2_1|r1[3]&r2[10]&add|r1[3]&r2[10]&sub|r1[3]&r2[10]&mul|r1[3]&r2[10]&act_func|r1[3]&r2[10]&act_func_2_1|r1[3]&r2[11]&add|r1[3]&r2[11]&sub|r1[3]&r2[11]&mul|r1[3]&r2[11]&act_func|r1[3]&r2[11]&act_func_2_1|r1[3]&r2[12]&add|r1[3]&r2[12]&sub|r1[3]&r2[12]&mul|r1[3]&r2[12]&act_func|r1[3]&r2[12]&act_func_2_1|r1[3]&r2[13]&sub|r1[3]&r2[13]&mul|r1[3]&r2[13]&act_func|r1[3]&r2[13]&act_func_2_1|r1[3]&r2[14]&sub|r1[3]&r2[14]&mul|r1[3]&r2[14]&act_func|r1[3]&r2[14]&act_func_2_1|r1[3]&r2[15]&sub|r1[3]&r2[15]&mul|r1[3]&r2[15]&act_func|r1[3]&r2[15]&act_func_2_1|r1[4]&r2[0]&add|r1[4]&r2[0]&sub|r1[4]&r2[0]&div|r1[4]&r2[0]&mul|r1[4]&r2[0]&pow|r1[4]&r2[0]&act_func|r1[4]&r2[0]&act_func_2_1|r1[4]&r2[1]&add|r1[4]&r2[1]&sub|r1[4]&r2[1]&div|r1[4]&r2[1]&mul|r1[4]&r2[1]&pow|r1[4]&r2[1]&act_func|r1[4]&r2[1]&act_func_2_1|r1[4]&r2[2]&add|r1[4]&r2[2]&sub|r1[4]&r2[2]&div|r1[4]&r2[2]&mul|r1[4]&r2[2]&act_func|r1[4]&r2[2]&act_func_2_1|r1[4]&r2[3]&add|r1[4]&r2[3]&sub|r1[4]&r2[3]&div|r1[4]&r2[3]&mul|r1[4]&r2[3]&pow|r1[4]&r2[3]&act_func|r1[4]&r2[3]&act_func_2_1|r1[4]&r2[4]&add|r1[4]&r2[4]&sub|r1[4]&r2[4]&mul|r1[4]&r2[4]&pow|r1[4]&r2[4]&act_func|r1[4]&r2[4]&act_func_2_1|r1[4]&r2[5]&add|r1[4]&r2[5]&sub|r1[4]&r2[5]&mul|r1[4]&r2[5]&pow|r1[4]&r2[5]&act_func|r1[4]&r2[5]&act_func_2_1|r1[4]&r2[6]&add|r1[4]&r2[6]&sub|r1[4]&r2[6]&mul|r1[4]&r2[6]&pow|r1[4]&r2[6]&act_func|r1[4]&r2[6]&act_func_2_1|r1[4]&r2[7]&add|r1[4]&r2[7]&sub|r1[4]&r2[7]&mul|r1[4]&r2[7]&pow|r1[4]&r2[7]&act_func|r1[4]&r2[7]&act_func_2_1|r1[4]&r2[8]&add|r1[4]&r2[8]&sub|r1[4]&r2[8]&mul|r1[4]&r2[8]&pow|r1[4]&r2[8]&act_func|r1[4]&r2[8]&act_func_2_1|r1[4]&r2[9]&add|r1[4]&r2[9]&sub|r1[4]&r2[9]&mul|r1[4]&r2[9]&pow|r1[4]&r2[9]&act_func|r1[4]&r2[9]&act_func_2_1|r1[4]&r2[10]&add|r1[4]&r2[10]&sub|r1[4]&r2[10]&mul|r1[4]&r2[10]&pow|r1[4]&r2[10]&act_func|r1[4]&r2[10]&act_func_2_1|r1[4]&r2[11]&add|r1[4]&r2[11]&sub|r1[4]&r2[11]&mul|r1[4]&r2[11]&pow|r1[4]&r2[11]&act_func|r1[4]&r2[11]&act_func_2_1|r1[4]&r2[12]&sub|r1[4]&r2[12]&mul|r1[4]&r2[12]&pow|r1[4]&r2[12]&act_func|r1[4]&r2[12]&act_func_2_1|r1[4]&r2[13]&sub|r1[4]&r2[13]&mul|r1[4]&r2[13]&pow|r1[4]&r2[13]&act_func|r1[4]&r2[13]&act_func_2_1|r1[4]&r2[14]&sub|r1[4]&r2[14]&mul|r1[4]&r2[14]&pow|r1[4]&r2[14]&act_func|r1[4]&r2[14]&act_func_2_1|r1[4]&r2[15]&sub|r1[4]&r2[15]&mul|r1[4]&r2[15]&pow|r1[4]&r2[15]&act_func|r1[4]&r2[15]&act_func_2_1|r1[5]&r2[0]&add|r1[5]&r2[0]&sub|r1[5]&r2[0]&div|r1[5]&r2[0]&mul|r1[5]&r2[0]&pow|r1[5]&r2[0]&act_func|r1[5]&r2[0]&act_func_2_1|r1[5]&r2[1]&add|r1[5]&r2[1]&sub|r1[5]&r2[1]&div|r1[5]&r2[1]&mul|r1[5]&r2[1]&pow|r1[5]&r2[1]&act_func|r1[5]&r2[1]&act_func_2_1|r1[5]&r2[2]&add|r1[5]&r2[2]&sub|r1[5]&r2[2]&div|r1[5]&r2[2]&mul|r1[5]&r2[2]&act_func|r1[5]&r2[2]&act_func_2_1|r1[5]&r2[3]&add|r1[5]&r2[3]&sub|r1[5]&r2[3]&div|r1[5]&r2[3]&mul|r1[5]&r2[3]&act_func|r1[5]&r2[3]&act_func_2_1|r1[5]&r2[4]&add|r1[5]&r2[4]&sub|r1[5]&r2[4]&mul|r1[5]&r2[4]&act_func|r1[5]&r2[4]&act_func_2_1|r1[5]&r2[5]&add|r1[5]&r2[5]&sub|r1[5]&r2[5]&mul|r1[5]&r2[5]&act_func|r1[5]&r2[5]&act_func_2_1|r1[5]&r2[6]&add|r1[5]&r2[6]&sub|r1[5]&r2[6]&mul|r1[5]&r2[6]&pow|r1[5]&r2[6]&act_func|r1[5]&r2[6]&act_func_2_1|r1[5]&r2[7]&add|r1[5]&r2[7]&sub|r1[5]&r2[7]&mul|r1[5]&r2[7]&act_func|r1[5]&r2[7]&act_func_2_1|r1[5]&r2[8]&add|r1[5]&r2[8]&sub|r1[5]&r2[8]&mul|r1[5]&r2[8]&act_func|r1[5]&r2[8]&act_func_2_1|r1[5]&r2[9]&add|r1[5]&r2[9]&sub|r1[5]&r2[9]&mul|r1[5]&r2[9]&act_func|r1[5]&r2[9]&act_func_2_1|r1[5]&r2[10]&add|r1[5]&r2[10]&sub|r1[5]&r2[10]&mul|r1[5]&r2[10]&act_func|r1[5]&r2[10]&act_func_2_1|r1[5]&r2[11]&sub|r1[5]&r2[11]&mul|r1[5]&r2[11]&act_func|r1[5]&r2[11]&act_func_2_1|r1[5]&r2[12]&sub|r1[5]&r2[12]&mul|r1[5]&r2[12]&act_func|r1[5]&r2[12]&act_func_2_1|r1[5]&r2[13]&sub|r1[5]&r2[13]&div|r1[5]&r2[13]&mul|r1[5]&r2[13]&act_func|r1[5]&r2[13]&act_func_2_1|r1[5]&r2[14]&sub|r1[5]&r2[14]&div|r1[5]&r2[14]&mul|r1[5]&r2[14]&act_func|r1[5]&r2[14]&act_func_2_1|r1[5]&r2[15]&sub|r1[5]&r2[15]&div|r1[5]&r2[15]&mul|r1[5]&r2[15]&pow|r1[5]&r2[15]&act_func|r1[5]&r2[15]&act_func_2_1|r1[6]&r2[0]&add|r1[6]&r2[0]&sub|r1[6]&r2[0]&div|r1[6]&r2[0]&mul|r1[6]&r2[0]&pow|r1[6]&r2[0]&act_func|r1[6]&r2[0]&act_func_2_1|r1[6]&r2[1]&add|r1[6]&r2[1]&sub|r1[6]&r2[1]&div|r1[6]&r2[1]&mul|r1[6]&r2[1]&pow|r1[6]&r2[1]&act_func|r1[6]&r2[1]&act_func_2_1|r1[6]&r2[2]&add|r1[6]&r2[2]&sub|r1[6]&r2[2]&div|r1[6]&r2[2]&mul|r1[6]&r2[2]&act_func|r1[6]&r2[2]&act_func_2_1|r1[6]&r2[3]&add|r1[6]&r2[3]&sub|r1[6]&r2[3]&mul|r1[6]&r2[3]&act_func|r1[6]&r2[3]&act_func_2_1|r1[6]&r2[4]&add|r1[6]&r2[4]&sub|r1[6]&r2[4]&mul|r1[6]&r2[4]&act_func|r1[6]&r2[4]&act_func_2_1|r1[6]&r2[5]&add|r1[6]&r2[5]&sub|r1[6]&r2[5]&mul|r1[6]&r2[5]&act_func|r1[6]&r2[5]&act_func_2_1|r1[6]&r2[6]&add|r1[6]&r2[6]&sub|r1[6]&r2[6]&mul|r1[6]&r2[6]&pow|r1[6]&r2[6]&act_func|r1[6]&r2[6]&act_func_2_1|r1[6]&r2[7]&add|r1[6]&r2[7]&sub|r1[6]&r2[7]&mul|r1[6]&r2[7]&pow|r1[6]&r2[7]&act_func|r1[6]&r2[7]&act_func_2_1|r1[6]&r2[8]&add|r1[6]&r2[8]&sub|r1[6]&r2[8]&mul|r1[6]&r2[8]&pow|r1[6]&r2[8]&act_func|r1[6]&r2[8]&act_func_2_1|r1[6]&r2[9]&add|r1[6]&r2[9]&sub|r1[6]&r2[9]&mul|r1[6]&r2[9]&pow|r1[6]&r2[9]&act_func|r1[6]&r2[9]&act_func_2_1|r1[6]&r2[10]&sub|r1[6]&r2[10]&mul|r1[6]&r2[10]&pow|r1[6]&r2[10]&act_func|r1[6]&r2[10]&act_func_2_1|r1[6]&r2[11]&sub|r1[6]&r2[11]&div|r1[6]&r2[11]&mul|r1[6]&r2[11]&pow|r1[6]&r2[11]&act_func|r1[6]&r2[11]&act_func_2_1|r1[6]&r2[12]&sub|r1[6]&r2[12]&div|r1[6]&r2[12]&mul|r1[6]&r2[12]&pow|r1[6]&r2[12]&act_func|r1[6]&r2[12]&act_func_2_1|r1[6]&r2[13]&sub|r1[6]&r2[13]&div|r1[6]&r2[13]&mul|r1[6]&r2[13]&pow|r1[6]&r2[13]&act_func|r1[6]&r2[13]&act_func_2_1|r1[6]&r2[14]&sub|r1[6]&r2[14]&mul|r1[6]&r2[14]&pow|r1[6]&r2[14]&act_func|r1[6]&r2[14]&act_func_2_1|r1[6]&r2[15]&sub|r1[6]&r2[15]&mul|r1[6]&r2[15]&pow|r1[6]&r2[15]&act_func|r1[6]&r2[15]&act_func_2_1|r1[7]&r2[0]&add|r1[7]&r2[0]&sub|r1[7]&r2[0]&div|r1[7]&r2[0]&mul|r1[7]&r2[0]&pow|r1[7]&r2[0]&act_func|r1[7]&r2[0]&act_func_2_1|r1[7]&r2[1]&add|r1[7]&r2[1]&sub|r1[7]&r2[1]&div|r1[7]&r2[1]&mul|r1[7]&r2[1]&pow|r1[7]&r2[1]&act_func|r1[7]&r2[1]&act_func_2_1|r1[7]&r2[2]&add|r1[7]&r2[2]&sub|r1[7]&r2[2]&div|r1[7]&r2[2]&mul|r1[7]&r2[2]&act_func|r1[7]&r2[2]&act_func_2_1|r1[7]&r2[3]&add|r1[7]&r2[3]&sub|r1[7]&r2[3]&mul|r1[7]&r2[3]&act_func|r1[7]&r2[3]&act_func_2_1|r1[7]&r2[4]&add|r1[7]&r2[4]&sub|r1[7]&r2[4]&mul|r1[7]&r2[4]&act_func|r1[7]&r2[4]&act_func_2_1|r1[7]&r2[5]&add|r1[7]&r2[5]&sub|r1[7]&r2[5]&mul|r1[7]&r2[5]&act_func|r1[7]&r2[5]&act_func_2_1|r1[7]&r2[6]&add|r1[7]&r2[6]&sub|r1[7]&r2[6]&mul|r1[7]&r2[6]&act_func|r1[7]&r2[6]&act_func_2_1|r1[7]&r2[7]&add|r1[7]&r2[7]&sub|r1[7]&r2[7]&mul|r1[7]&r2[7]&act_func|r1[7]&r2[7]&act_func_2_1|r1[7]&r2[8]&add|r1[7]&r2[8]&sub|r1[7]&r2[8]&mul|r1[7]&r2[8]&pow|r1[7]&r2[8]&act_func|r1[7]&r2[8]&act_func_2_1|r1[7]&r2[9]&sub|r1[7]&r2[9]&mul|r1[7]&r2[9]&pow|r1[7]&r2[9]&act_func|r1[7]&r2[9]&act_func_2_1|r1[7]&r2[10]&sub|r1[7]&r2[10]&div|r1[7]&r2[10]&mul|r1[7]&r2[10]&act_func|r1[7]&r2[10]&act_func_2_1|r1[7]&r2[11]&sub|r1[7]&r2[11]&div|r1[7]&r2[11]&mul|r1[7]&r2[11]&act_func|r1[7]&r2[11]&act_func_2_1|r1[7]&r2[12]&sub|r1[7]&r2[12]&mul|r1[7]&r2[12]&act_func|r1[7]&r2[12]&act_func_2_1|r1[7]&r2[13]&sub|r1[7]&r2[13]&mul|r1[7]&r2[13]&act_func|r1[7]&r2[13]&act_func_2_1|r1[7]&r2[14]&sub|r1[7]&r2[14]&mul|r1[7]&r2[14]&act_func|r1[7]&r2[14]&act_func_2_1|r1[7]&r2[15]&sub|r1[7]&r2[15]&mul|r1[7]&r2[15]&act_func|r1[7]&r2[15]&act_func_2_1|r1[8]&r2[0]&add|r1[8]&r2[0]&sub|r1[8]&r2[0]&div|r1[8]&r2[0]&mul|r1[8]&r2[0]&pow|r1[8]&r2[0]&act_func|r1[8]&r2[0]&act_func_2_1|r1[8]&r2[1]&add|r1[8]&r2[1]&sub|r1[8]&r2[1]&div|r1[8]&r2[1]&mul|r1[8]&r2[1]&pow|r1[8]&r2[1]&act_func|r1[8]&r2[1]&act_func_2_1|r1[8]&r2[2]&add|r1[8]&r2[2]&sub|r1[8]&r2[2]&mul|r1[8]&r2[2]&pow|r1[8]&r2[2]&act_func|r1[8]&r2[2]&act_func_2_1|r1[8]&r2[3]&add|r1[8]&r2[3]&sub|r1[8]&r2[3]&mul|r1[8]&r2[3]&pow|r1[8]&r2[3]&act_func|r1[8]&r2[3]&act_func_2_1|r1[8]&r2[4]&add|r1[8]&r2[4]&sub|r1[8]&r2[4]&mul|r1[8]&r2[4]&pow|r1[8]&r2[4]&act_func|r1[8]&r2[4]&act_func_2_1|r1[8]&r2[5]&add|r1[8]&r2[5]&sub|r1[8]&r2[5]&mul|r1[8]&r2[5]&pow|r1[8]&r2[5]&act_func|r1[8]&r2[5]&act_func_2_1|r1[8]&r2[6]&add|r1[8]&r2[6]&sub|r1[8]&r2[6]&mul|r1[8]&r2[6]&pow|r1[8]&r2[6]&act_func|r1[8]&r2[6]&act_func_2_1|r1[8]&r2[7]&add|r1[8]&r2[7]&sub|r1[8]&r2[7]&mul|r1[8]&r2[7]&pow|r1[8]&r2[7]&act_func|r1[8]&r2[7]&act_func_2_1|r1[8]&r2[8]&sub|r1[8]&r2[8]&div|r1[8]&r2[8]&mul|r1[8]&r2[8]&pow|r1[8]&r2[8]&act_func|r1[8]&r2[8]&act_func_2_1|r1[8]&r2[9]&sub|r1[8]&r2[9]&div|r1[8]&r2[9]&mul|r1[8]&r2[9]&pow|r1[8]&r2[9]&act_func|r1[8]&r2[9]&act_func_2_1|r1[8]&r2[10]&sub|r1[8]&r2[10]&mul|r1[8]&r2[10]&pow|r1[8]&r2[10]&act_func|r1[8]&r2[10]&act_func_2_1|r1[8]&r2[11]&sub|r1[8]&r2[11]&mul|r1[8]&r2[11]&pow|r1[8]&r2[11]&act_func|r1[8]&r2[11]&act_func_2_1|r1[8]&r2[12]&sub|r1[8]&r2[12]&mul|r1[8]&r2[12]&pow|r1[8]&r2[12]&act_func|r1[8]&r2[12]&act_func_2_1|r1[8]&r2[13]&sub|r1[8]&r2[13]&mul|r1[8]&r2[13]&pow|r1[8]&r2[13]&act_func|r1[8]&r2[13]&act_func_2_1|r1[8]&r2[14]&sub|r1[8]&r2[14]&mul|r1[8]&r2[14]&pow|r1[8]&r2[14]&act_func|r1[8]&r2[14]&act_func_2_1|r1[8]&r2[15]&sub|r1[8]&r2[15]&mul|r1[8]&r2[15]&pow|r1[8]&r2[15]&act_func|r1[8]&r2[15]&act_func_2_1|r1[9]&r2[0]&add|r1[9]&r2[0]&sub|r1[9]&r2[0]&div|r1[9]&r2[0]&mul|r1[9]&r2[0]&pow|r1[9]&r2[0]&act_func|r1[9]&r2[0]&act_func_2_1|r1[9]&r2[1]&add|r1[9]&r2[1]&sub|r1[9]&r2[1]&div|r1[9]&r2[1]&mul|r1[9]&r2[1]&pow|r1[9]&r2[1]&act_func|r1[9]&r2[1]&act_func_2_1|r1[9]&r2[2]&add|r1[9]&r2[2]&sub|r1[9]&r2[2]&mul|r1[9]&r2[2]&act_func|r1[9]&r2[2]&act_func_2_1|r1[9]&r2[3]&add|r1[9]&r2[3]&sub|r1[9]&r2[3]&mul|r1[9]&r2[3]&act_func|r1[9]&r2[3]&act_func_2_1|r1[9]&r2[4]&add|r1[9]&r2[4]&sub|r1[9]&r2[4]&mul|r1[9]&r2[4]&act_func|r1[9]&r2[4]&act_func_2_1|r1[9]&r2[5]&add|r1[9]&r2[5]&sub|r1[9]&r2[5]&mul|r1[9]&r2[5]&act_func|r1[9]&r2[5]&act_func_2_1|r1[9]&r2[6]&add|r1[9]&r2[6]&sub|r1[9]&r2[6]&mul|r1[9]&r2[6]&act_func|r1[9]&r2[6]&act_func_2_1|r1[9]&r2[7]&sub|r1[9]&r2[7]&mul|r1[9]&r2[7]&act_func|r1[9]&r2[7]&act_func_2_1|r1[9]&r2[8]&sub|r1[9]&r2[8]&div|r1[9]&r2[8]&mul|r1[9]&r2[8]&pow|r1[9]&r2[8]&act_func|r1[9]&r2[8]&act_func_2_1|r1[9]&r2[9]&sub|r1[9]&r2[9]&mul|r1[9]&r2[9]&pow|r1[9]&r2[9]&act_func|r1[9]&r2[9]&act_func_2_1|r1[9]&r2[10]&sub|r1[9]&r2[10]&mul|r1[9]&r2[10]&act_func|r1[9]&r2[10]&act_func_2_1|r1[9]&r2[11]&sub|r1[9]&r2[11]&mul|r1[9]&r2[11]&act_func|r1[9]&r2[11]&act_func_2_1|r1[9]&r2[12]&sub|r1[9]&r2[12]&mul|r1[9]&r2[12]&act_func|r1[9]&r2[12]&act_func_2_1|r1[9]&r2[13]&sub|r1[9]&r2[13]&mul|r1[9]&r2[13]&act_func|r1[9]&r2[13]&act_func_2_1|r1[9]&r2[14]&sub|r1[9]&r2[14]&mul|r1[9]&r2[14]&act_func|r1[9]&r2[14]&act_func_2_1|r1[9]&r2[15]&sub|r1[9]&r2[15]&div|r1[9]&r2[15]&mul|r1[9]&r2[15]&act_func|r1[9]&r2[15]&act_func_2_1|r1[10]&r2[0]&add|r1[10]&r2[0]&sub|r1[10]&r2[0]&div|r1[10]&r2[0]&mul|r1[10]&r2[0]&pow|r1[10]&r2[0]&act_func|r1[10]&r2[0]&act_func_2_1|r1[10]&r2[1]&add|r1[10]&r2[1]&sub|r1[10]&r2[1]&div|r1[10]&r2[1]&mul|r1[10]&r2[1]&pow|r1[10]&r2[1]&act_func|r1[10]&r2[1]&act_func_2_1|r1[10]&r2[2]&add|r1[10]&r2[2]&sub|r1[10]&r2[2]&mul|r1[10]&r2[2]&act_func|r1[10]&r2[2]&act_func_2_1|r1[10]&r2[3]&add|r1[10]&r2[3]&sub|r1[10]&r2[3]&mul|r1[10]&r2[3]&act_func|r1[10]&r2[3]&act_func_2_1|r1[10]&r2[4]&add|r1[10]&r2[4]&sub|r1[10]&r2[4]&mul|r1[10]&r2[4]&act_func|r1[10]&r2[4]&act_func_2_1|r1[10]&r2[5]&add|r1[10]&r2[5]&sub|r1[10]&r2[5]&mul|r1[10]&r2[5]&act_func|r1[10]&r2[5]&act_func_2_1|r1[10]&r2[6]&sub|r1[10]&r2[6]&mul|r1[10]&r2[6]&pow|r1[10]&r2[6]&act_func|r1[10]&r2[6]&act_func_2_1|r1[10]&r2[7]&sub|r1[10]&r2[7]&div|r1[10]&r2[7]&mul|r1[10]&r2[7]&pow|r1[10]&r2[7]&act_func|r1[10]&r2[7]&act_func_2_1|r1[10]&r2[8]&sub|r1[10]&r2[8]&mul|r1[10]&r2[8]&pow|r1[10]&r2[8]&act_func|r1[10]&r2[8]&act_func_2_1|r1[10]&r2[9]&sub|r1[10]&r2[9]&mul|r1[10]&r2[9]&pow|r1[10]&r2[9]&act_func|r1[10]&r2[9]&act_func_2_1|r1[10]&r2[10]&sub|r1[10]&r2[10]&mul|r1[10]&r2[10]&pow|r1[10]&r2[10]&act_func|r1[10]&r2[10]&act_func_2_1|r1[10]&r2[11]&sub|r1[10]&r2[11]&mul|r1[10]&r2[11]&pow|r1[10]&r2[11]&act_func|r1[10]&r2[11]&act_func_2_1|r1[10]&r2[12]&sub|r1[10]&r2[12]&mul|r1[10]&r2[12]&pow|r1[10]&r2[12]&act_func|r1[10]&r2[12]&act_func_2_1|r1[10]&r2[13]&sub|r1[10]&r2[13]&div|r1[10]&r2[13]&mul|r1[10]&r2[13]&pow|r1[10]&r2[13]&act_func|r1[10]&r2[13]&act_func_2_1|r1[10]&r2[14]&sub|r1[10]&r2[14]&div|r1[10]&r2[14]&mul|r1[10]&r2[14]&pow|r1[10]&r2[14]&act_func|r1[10]&r2[14]&act_func_2_1|r1[10]&r2[15]&sub|r1[10]&r2[15]&mul|r1[10]&r2[15]&pow|r1[10]&r2[15]&act_func|r1[10]&r2[15]&act_func_2_1|r1[11]&r2[0]&add|r1[11]&r2[0]&sub|r1[11]&r2[0]&div|r1[11]&r2[0]&mul|r1[11]&r2[0]&pow|r1[11]&r2[0]&act_func|r1[11]&r2[0]&act_func_2_1|r1[11]&r2[1]&add|r1[11]&r2[1]&sub|r1[11]&r2[1]&div|r1[11]&r2[1]&mul|r1[11]&r2[1]&pow|r1[11]&r2[1]&act_func|r1[11]&r2[1]&act_func_2_1|r1[11]&r2[2]&add|r1[11]&r2[2]&sub|r1[11]&r2[2]&mul|r1[11]&r2[2]&act_func|r1[11]&r2[2]&act_func_2_1|r1[11]&r2[3]&add|r1[11]&r2[3]&sub|r1[11]&r2[3]&mul|r1[11]&r2[3]&act_func|r1[11]&r2[3]&act_func_2_1|r1[11]&r2[4]&add|r1[11]&r2[4]&sub|r1[11]&r2[4]&mul|r1[11]&r2[4]&act_func|r1[11]&r2[4]&act_func_2_1|r1[11]&r2[5]&sub|r1[11]&r2[5]&mul|r1[11]&r2[5]&act_func|r1[11]&r2[5]&act_func_2_1|r1[11]&r2[6]&sub|r1[11]&r2[6]&div|r1[11]&r2[6]&mul|r1[11]&r2[6]&act_func|r1[11]&r2[6]&act_func_2_1|r1[11]&r2[7]&sub|r1[11]&r2[7]&div|r1[11]&r2[7]&mul|r1[11]&r2[7]&pow|r1[11]&r2[7]&act_func|r1[11]&r2[7]&act_func_2_1|r1[11]&r2[8]&sub|r1[11]&r2[8]&mul|r1[11]&r2[8]&act_func|r1[11]&r2[8]&act_func_2_1|r1[11]&r2[9]&sub|r1[11]&r2[9]&mul|r1[11]&r2[9]&act_func|r1[11]&r2[9]&act_func_2_1|r1[11]&r2[10]&sub|r1[11]&r2[10]&mul|r1[11]&r2[10]&act_func|r1[11]&r2[10]&act_func_2_1|r1[11]&r2[11]&sub|r1[11]&r2[11]&mul|r1[11]&r2[11]&act_func|r1[11]&r2[11]&act_func_2_1|r1[11]&r2[12]&sub|r1[11]&r2[12]&div|r1[11]&r2[12]&mul|r1[11]&r2[12]&act_func|r1[11]&r2[12]&act_func_2_1|r1[11]&r2[13]&sub|r1[11]&r2[13]&div|r1[11]&r2[13]&mul|r1[11]&r2[13]&act_func|r1[11]&r2[13]&act_func_2_1|r1[11]&r2[14]&sub|r1[11]&r2[14]&mul|r1[11]&r2[14]&pow|r1[11]&r2[14]&act_func|r1[11]&r2[14]&act_func_2_1|r1[11]&r2[15]&sub|r1[11]&r2[15]&mul|r1[11]&r2[15]&act_func|r1[11]&r2[15]&act_func_2_1|r1[12]&r2[0]&add|r1[12]&r2[0]&sub|r1[12]&r2[0]&div|r1[12]&r2[0]&mul|r1[12]&r2[0]&pow|r1[12]&r2[0]&act_func|r1[12]&r2[0]&act_func_2_1|r1[12]&r2[1]&add|r1[12]&r2[1]&sub|r1[12]&r2[1]&div|r1[12]&r2[1]&mul|r1[12]&r2[1]&pow|r1[12]&r2[1]&act_func|r1[12]&r2[1]&act_func_2_1|r1[12]&r2[2]&add|r1[12]&r2[2]&sub|r1[12]&r2[2]&mul|r1[12]&r2[2]&act_func|r1[12]&r2[2]&act_func_2_1|r1[12]&r2[3]&add|r1[12]&r2[3]&sub|r1[12]&r2[3]&mul|r1[12]&r2[3]&pow|r1[12]&r2[3]&act_func|r1[12]&r2[3]&act_func_2_1|r1[12]&r2[4]&sub|r1[12]&r2[4]&mul|r1[12]&r2[4]&pow|r1[12]&r2[4]&act_func|r1[12]&r2[4]&act_func_2_1|r1[12]&r2[5]&sub|r1[12]&r2[5]&mul|r1[12]&r2[5]&pow|r1[12]&r2[5]&act_func|r1[12]&r2[5]&act_func_2_1|r1[12]&r2[6]&sub|r1[12]&r2[6]&div|r1[12]&r2[6]&mul|r1[12]&r2[6]&pow|r1[12]&r2[6]&act_func|r1[12]&r2[6]&act_func_2_1|r1[12]&r2[7]&sub|r1[12]&r2[7]&mul|r1[12]&r2[7]&pow|r1[12]&r2[7]&act_func|r1[12]&r2[7]&act_func_2_1|r1[12]&r2[8]&sub|r1[12]&r2[8]&mul|r1[12]&r2[8]&pow|r1[12]&r2[8]&act_func|r1[12]&r2[8]&act_func_2_1|r1[12]&r2[9]&sub|r1[12]&r2[9]&mul|r1[12]&r2[9]&pow|r1[12]&r2[9]&act_func|r1[12]&r2[9]&act_func_2_1|r1[12]&r2[10]&sub|r1[12]&r2[10]&mul|r1[12]&r2[10]&pow|r1[12]&r2[10]&act_func|r1[12]&r2[10]&act_func_2_1|r1[12]&r2[11]&sub|r1[12]&r2[11]&div|r1[12]&r2[11]&mul|r1[12]&r2[11]&pow|r1[12]&r2[11]&act_func|r1[12]&r2[11]&act_func_2_1|r1[12]&r2[12]&sub|r1[12]&r2[12]&mul|r1[12]&r2[12]&pow|r1[12]&r2[12]&act_func|r1[12]&r2[12]&act_func_2_1|r1[12]&r2[13]&sub|r1[12]&r2[13]&mul|r1[12]&r2[13]&pow|r1[12]&r2[13]&act_func|r1[12]&r2[13]&act_func_2_1|r1[12]&r2[14]&sub|r1[12]&r2[14]&mul|r1[12]&r2[14]&pow|r1[12]&r2[14]&act_func|r1[12]&r2[14]&act_func_2_1|r1[12]&r2[15]&sub|r1[12]&r2[15]&mul|r1[12]&r2[15]&pow|r1[12]&r2[15]&act_func|r1[12]&r2[15]&act_func_2_1|r1[13]&r2[0]&add|r1[13]&r2[0]&sub|r1[13]&r2[0]&div|r1[13]&r2[0]&mul|r1[13]&r2[0]&pow|r1[13]&r2[0]&act_func|r1[13]&r2[0]&act_func_2_1|r1[13]&r2[1]&add|r1[13]&r2[1]&sub|r1[13]&r2[1]&div|r1[13]&r2[1]&mul|r1[13]&r2[1]&pow|r1[13]&r2[1]&act_func|r1[13]&r2[1]&act_func_2_1|r1[13]&r2[2]&add|r1[13]&r2[2]&sub|r1[13]&r2[2]&mul|r1[13]&r2[2]&act_func|r1[13]&r2[2]&act_func_2_1|r1[13]&r2[3]&sub|r1[13]&r2[3]&mul|r1[13]&r2[3]&act_func|r1[13]&r2[3]&act_func_2_1|r1[13]&r2[4]&sub|r1[13]&r2[4]&mul|r1[13]&r2[4]&act_func|r1[13]&r2[4]&act_func_2_1|r1[13]&r2[5]&sub|r1[13]&r2[5]&div|r1[13]&r2[5]&mul|r1[13]&r2[5]&act_func|r1[13]&r2[5]&act_func_2_1|r1[13]&r2[6]&sub|r1[13]&r2[6]&div|r1[13]&r2[6]&mul|r1[13]&r2[6]&act_func|r1[13]&r2[6]&act_func_2_1|r1[13]&r2[7]&sub|r1[13]&r2[7]&mul|r1[13]&r2[7]&act_func|r1[13]&r2[7]&act_func_2_1|r1[13]&r2[8]&sub|r1[13]&r2[8]&mul|r1[13]&r2[8]&act_func|r1[13]&r2[8]&act_func_2_1|r1[13]&r2[9]&sub|r1[13]&r2[9]&mul|r1[13]&r2[9]&act_func|r1[13]&r2[9]&act_func_2_1|r1[13]&r2[10]&sub|r1[13]&r2[10]&div|r1[13]&r2[10]&mul|r1[13]&r2[10]&pow|r1[13]&r2[10]&act_func|r1[13]&r2[10]&act_func_2_1|r1[13]&r2[11]&sub|r1[13]&r2[11]&div|r1[13]&r2[11]&mul|r1[13]&r2[11]&act_func|r1[13]&r2[11]&act_func_2_1|r1[13]&r2[12]&sub|r1[13]&r2[12]&mul|r1[13]&r2[12]&act_func|r1[13]&r2[12]&act_func_2_1|r1[13]&r2[13]&sub|r1[13]&r2[13]&mul|r1[13]&r2[13]&act_func|r1[13]&r2[13]&act_func_2_1|r1[13]&r2[14]&sub|r1[13]&r2[14]&mul|r1[13]&r2[14]&act_func|r1[13]&r2[14]&act_func_2_1|r1[13]&r2[15]&sub|r1[13]&r2[15]&div|r1[13]&r2[15]&mul|r1[13]&r2[15]&pow|r1[13]&r2[15]&act_func|r1[13]&r2[15]&act_func_2_1|r1[14]&r2[0]&add|r1[14]&r2[0]&sub|r1[14]&r2[0]&div|r1[14]&r2[0]&mul|r1[14]&r2[0]&pow|r1[14]&r2[0]&act_func|r1[14]&r2[0]&act_func_2_1|r1[14]&r2[1]&add|r1[14]&r2[1]&sub|r1[14]&r2[1]&div|r1[14]&r2[1]&mul|r1[14]&r2[1]&pow|r1[14]&r2[1]&act_func|r1[14]&r2[1]&act_func_2_1|r1[14]&r2[2]&sub|r1[14]&r2[2]&mul|r1[14]&r2[2]&pow|r1[14]&r2[2]&act_func|r1[14]&r2[2]&act_func_2_1|r1[14]&r2[3]&sub|r1[14]&r2[3]&mul|r1[14]&r2[3]&act_func|r1[14]&r2[3]&act_func_2_1|r1[14]&r2[4]&sub|r1[14]&r2[4]&mul|r1[14]&r2[4]&act_func|r1[14]&r2[4]&act_func_2_1|r1[14]&r2[5]&sub|r1[14]&r2[5]&div|r1[14]&r2[5]&mul|r1[14]&r2[5]&act_func|r1[14]&r2[5]&act_func_2_1|r1[14]&r2[6]&sub|r1[14]&r2[6]&mul|r1[14]&r2[6]&pow|r1[14]&r2[6]&act_func|r1[14]&r2[6]&act_func_2_1|r1[14]&r2[7]&sub|r1[14]&r2[7]&mul|r1[14]&r2[7]&pow|r1[14]&r2[7]&act_func|r1[14]&r2[7]&act_func_2_1|r1[14]&r2[8]&sub|r1[14]&r2[8]&mul|r1[14]&r2[8]&pow|r1[14]&r2[8]&act_func|r1[14]&r2[8]&act_func_2_1|r1[14]&r2[9]&sub|r1[14]&r2[9]&mul|r1[14]&r2[9]&pow|r1[14]&r2[9]&act_func|r1[14]&r2[9]&act_func_2_1|r1[14]&r2[10]&sub|r1[14]&r2[10]&div|r1[14]&r2[10]&mul|r1[14]&r2[10]&pow|r1[14]&r2[10]&act_func|r1[14]&r2[10]&act_func_2_1|r1[14]&r2[11]&sub|r1[14]&r2[11]&mul|r1[14]&r2[11]&pow|r1[14]&r2[11]&act_func|r1[14]&r2[11]&act_func_2_1|r1[14]&r2[12]&sub|r1[14]&r2[12]&mul|r1[14]&r2[12]&pow|r1[14]&r2[12]&act_func|r1[14]&r2[12]&act_func_2_1|r1[14]&r2[13]&sub|r1[14]&r2[13]&mul|r1[14]&r2[13]&pow|r1[14]&r2[13]&act_func|r1[14]&r2[13]&act_func_2_1|r1[14]&r2[14]&sub|r1[14]&r2[14]&div|r1[14]&r2[14]&mul|r1[14]&r2[14]&pow|r1[14]&r2[14]&act_func|r1[14]&r2[14]&act_func_2_1|r1[14]&r2[15]&sub|r1[14]&r2[15]&mul|r1[14]&r2[15]&pow|r1[14]&r2[15]&act_func|r1[14]&r2[15]&act_func_2_1|r1[15]&r2[0]&add|r1[15]&r2[0]&sub|r1[15]&r2[0]&div|r1[15]&r2[0]&mul|r1[15]&r2[0]&pow|r1[15]&r2[0]&act_func|r1[15]&r2[0]&act_func_2_1|r1[15]&r2[1]&sub|r1[15]&r2[1]&div|r1[15]&r2[1]&mul|r1[15]&r2[1]&pow|r1[15]&r2[1]&act_func|r1[15]&r2[1]&act_func_2_1|r1[15]&r2[2]&sub|r1[15]&r2[2]&mul|r1[15]&r2[2]&act_func|r1[15]&r2[2]&act_func_2_1|r1[15]&r2[3]&sub|r1[15]&r2[3]&mul|r1[15]&r2[3]&act_func|r1[15]&r2[3]&act_func_2_1|r1[15]&r2[4]&sub|r1[15]&r2[4]&mul|r1[15]&r2[4]&pow|r1[15]&r2[4]&act_func|r1[15]&r2[4]&act_func_2_1|r1[15]&r2[5]&sub|r1[15]&r2[5]&div|r1[15]&r2[5]&mul|r1[15]&r2[5]&pow|r1[15]&r2[5]&act_func|r1[15]&r2[5]&act_func_2_1|r1[15]&r2[6]&sub|r1[15]&r2[6]&mul|r1[15]&r2[6]&act_func|r1[15]&r2[6]&act_func_2_1|r1[15]&r2[7]&sub|r1[15]&r2[7]&mul|r1[15]&r2[7]&act_func|r1[15]&r2[7]&act_func_2_1|r1[15]&r2[8]&sub|r1[15]&r2[8]&mul|r1[15]&r2[8]&pow|r1[15]&r2[8]&act_func|r1[15]&r2[8]&act_func_2_1|r1[15]&r2[9]&sub|r1[15]&r2[9]&div|r1[15]&r2[9]&mul|r1[15]&r2[9]&pow|r1[15]&r2[9]&act_func|r1[15]&r2[9]&act_func_2_1|r1[15]&r2[10]&sub|r1[15]&r2[10]&mul|r1[15]&r2[10]&act_func|r1[15]&r2[10]&act_func_2_1|r1[15]&r2[11]&sub|r1[15]&r2[11]&mul|r1[15]&r2[11]&act_func|r1[15]&r2[11]&act_func_2_1|r1[15]&r2[12]&sub|r1[15]&r2[12]&mul|r1[15]&r2[12]&pow|r1[15]&r2[12]&act_func|r1[15]&r2[12]&act_func_2_1|r1[15]&r2[13]&sub|r1[15]&r2[13]&div|r1[15]&r2[13]&mul|r1[15]&r2[13]&pow|r1[15]&r2[13]&act_func|r1[15]&r2[13]&act_func_2_1|r1[15]&r2[14]&sub|r1[15]&r2[14]&mul|r1[15]&r2[14]&act_func|r1[15]&r2[14]&act_func_2_1|r1[15]&r2[15]&sub|r1[15]&r2[15]&mul|r1[15]&r2[15]&pow|r1[15]&r2[15]&act_func|r1[15]&r2[15]&act_func_2_1,
r1[0]&r2[15]&add|r1[1]&r2[14]&add|r1[1]&r2[15]&div|r1[2]&r2[13]&add|r1[3]&r2[5]&div|r1[3]&r2[12]&add|r1[4]&r2[11]&add|r1[5]&r2[3]&div|r1[5]&r2[10]&add|r1[6]&r2[9]&add|r1[7]&r2[8]&add|r1[7]&r2[9]&div|r1[8]&r2[7]&add|r1[9]&r2[6]&add|r1[9]&r2[7]&div|r1[10]&r2[5]&add|r1[11]&r2[4]&add|r1[11]&r2[13]&div|r1[12]&r2[3]&add|r1[13]&r2[2]&add|r1[13]&r2[11]&div|r1[14]&r2[1]&add|r1[15]&r2[0]&add|r1[15]&r2[0]&sub|r1[15]&r2[0]&mul|r1[15]&r2[1]&div|r1[15]&r2[1]&pow|r1[15]&r2[3]&pow|r1[15]&r2[5]&pow|r1[15]&r2[7]&pow|r1[15]&r2[9]&pow|r1[15]&r2[11]&pow|r1[15]&r2[13]&pow,
r1[0]&r2[14]&add|r1[1]&r2[13]&add|r1[1]&r2[14]&div|r1[2]&r2[7]&div|r1[2]&r2[12]&add|r1[2]&r2[15]&div|r1[3]&r2[10]&div|r1[3]&r2[11]&add|r1[4]&r2[10]&add|r1[5]&r2[6]&div|r1[5]&r2[9]&add|r1[6]&r2[5]&div|r1[6]&r2[8]&add|r1[6]&r2[13]&div|r1[7]&r2[2]&div|r1[7]&r2[7]&add|r1[8]&r2[6]&add|r1[9]&r2[5]&add|r1[9]&r2[14]&div|r1[10]&r2[3]&div|r1[10]&r2[4]&add|r1[10]&r2[11]&div|r1[11]&r2[3]&add|r1[11]&r2[10]&div|r1[12]&r2[2]&add|r1[13]&r2[1]&add|r1[13]&r2[6]&div|r1[14]&r2[0]&add|r1[14]&r2[0]&sub|r1[14]&r2[0]&mul|r1[14]&r2[1]&div|r1[14]&r2[1]&pow|r1[14]&r2[9]&div|r1[15]&r2[1]&sub|r1[15]&r2[2]&div|r1[15]&r2[15]&add,
r1[0]&r2[13]&add|r1[1]&r2[12]&add|r1[1]&r2[13]&div|r1[2]&r2[11]&add|r1[3]&r2[10]&add|r1[3]&r2[15]&div|r1[4]&r2[9]&add|r1[5]&r2[3]&pow|r1[5]&r2[7]&pow|r1[5]&r2[8]&add|r1[5]&r2[9]&div|r1[5]&r2[11]&pow|r1[5]&r2[15]&pow|r1[6]&r2[7]&add|r1[7]&r2[6]&add|r1[7]&r2[11]&div|r1[8]&r2[5]&add|r1[9]&r2[4]&add|r1[9]&r2[5]&div|r1[10]&r2[3]&add|r1[11]&r2[2]&add|r1[11]&r2[7]&div|r1[12]&r2[1]&add|r1[13]&r2[0]&add|r1[13]&r2[0]&sub|r1[13]&r2[0]&mul|r1[13]&r2[1]&div|r1[13]&r2[1]&pow|r1[13]&r2[5]&pow|r1[13]&r2[9]&pow|r1[13]&r2[13]&pow|r1[14]&r2[1]&sub|r1[14]&r2[15]&add|r1[15]&r2[2]&sub|r1[15]&r2[3]&div|r1[15]&r2[14]&add,
r1[0]&r2[12]&add|r1[1]&r2[11]&add|r1[1]&r2[12]&div|r1[2]&r2[6]&div|r1[2]&r2[10]&add|r1[2]&r2[14]&div|r1[3]&r2[4]&div|r1[3]&r2[9]&add|r1[4]&r2[3]&div|r1[4]&r2[7]&div|r1[4]&r2[8]&add|r1[4]&r2[11]&div|r1[4]&r2[15]&div|r1[5]&r2[7]&add|r1[5]&r2[12]&div|r1[6]&r2[2]&div|r1[6]&r2[6]&add|r1[6]&r2[10]&div|r1[7]&r2[4]&div|r1[7]&r2[5]&add|r1[8]&r2[4]&add|r1[9]&r2[3]&add|r1[9]&r2[12]&div|r1[10]&r2[2]&add|r1[10]&r2[6]&div|r1[10]&r2[14]&div|r1[11]&r2[1]&add|r1[11]&r2[4]&div|r1[12]&r2[0]&add|r1[12]&r2[0]&sub|r1[12]&r2[0]&mul|r1[12]&r2[1]&div|r1[12]&r2[1]&pow|r1[12]&r2[5]&div|r1[12]&r2[9]&div|r1[12]&r2[13]&div|r1[13]&r2[1]&sub|r1[13]&r2[12]&div|r1[13]&r2[15]&add|r1[14]&r2[2]&sub|r1[14]&r2[2]&div|r1[14]&r2[10]&div|r1[14]&r2[14]&add|r1[15]&r2[3]&sub|r1[15]&r2[4]&div|r1[15]&r2[13]&add,
r1[0]&r2[11]&add|r1[1]&r2[10]&add|r1[1]&r2[11]&div|r1[2]&r2[9]&add|r1[3]&r2[3]&pow|r1[3]&r2[7]&pow|r1[3]&r2[8]&add|r1[3]&r2[9]&div|r1[3]&r2[11]&pow|r1[3]&r2[15]&pow|r1[4]&r2[7]&add|r1[5]&r2[6]&add|r1[5]&r2[15]&div|r1[6]&r2[5]&add|r1[7]&r2[4]&add|r1[7]&r2[13]&div|r1[8]&r2[3]&add|r1[9]&r2[2]&add|r1[9]&r2[3]&div|r1[10]&r2[1]&add|r1[11]&r2[0]&add|r1[11]&r2[0]&sub|r1[11]&r2[0]&mul|r1[11]&r2[1]&div|r1[11]&r2[1]&pow|r1[11]&r2[5]&pow|r1[11]&r2[9]&pow|r1[11]&r2[13]&pow|r1[12]&r2[1]&sub|r1[12]&r2[15]&add|r1[13]&r2[2]&sub|r1[13]&r2[7]&div|r1[13]&r2[14]&add|r1[14]&r2[3]&sub|r1[14]&r2[13]&add|r1[15]&r2[4]&sub|r1[15]&r2[5]&div|r1[15]&r2[12]&add,
r1[0]&r2[10]&add|r1[1]&r2[9]&add|r1[1]&r2[10]&div|r1[2]&r2[5]&div|r1[2]&r2[8]&add|r1[2]&r2[13]&div|r1[3]&r2[7]&add|r1[3]&r2[14]&div|r1[4]&r2[6]&add|r1[5]&r2[2]&div|r1[5]&r2[5]&add|r1[6]&r2[4]&add|r1[6]&r2[7]&div|r1[6]&r2[15]&div|r1[7]&r2[3]&add|r1[7]&r2[6]&div|r1[8]&r2[2]&add|r1[9]&r2[1]&add|r1[9]&r2[10]&div|r1[10]&r2[0]&add|r1[10]&r2[0]&sub|r1[10]&r2[0]&mul|r1[10]&r2[1]&div|r1[10]&r2[1]&pow|r1[10]&r2[9]&div|r1[11]&r2[1]&sub|r1[11]&r2[14]&div|r1[11]&r2[15]&add|r1[12]&r2[2]&sub|r1[12]&r2[14]&add|r1[13]&r2[2]&div|r1[13]&r2[3]&sub|r1[13]&r2[13]&add|r1[14]&r2[3]&div|r1[14]&r2[4]&sub|r1[14]&r2[11]&div|r1[14]&r2[12]&add|r1[15]&r2[5]&sub|r1[15]&r2[6]&div|r1[15]&r2[11]&add,
r1[0]&r2[9]&add|r1[1]&r2[8]&add|r1[1]&r2[9]&div|r1[2]&r2[7]&add|r1[3]&r2[2]&pow|r1[3]&r2[3]&div|r1[3]&r2[6]&add|r1[3]&r2[6]&pow|r1[3]&r2[10]&pow|r1[3]&r2[14]&pow|r1[4]&r2[5]&add|r1[5]&r2[2]&pow|r1[5]&r2[4]&add|r1[5]&r2[5]&div|r1[5]&r2[6]&pow|r1[5]&r2[10]&pow|r1[5]&r2[14]&pow|r1[6]&r2[3]&add|r1[7]&r2[2]&add|r1[7]&r2[15]&div|r1[8]&r2[1]&add|r1[9]&r2[0]&add|r1[9]&r2[0]&sub|r1[9]&r2[0]&mul|r1[9]&r2[1]&div|r1[9]&r2[1]&pow|r1[9]&r2[3]&pow|r1[9]&r2[5]&pow|r1[9]&r2[7]&pow|r1[9]&r2[9]&pow|r1[9]&r2[11]&pow|r1[9]&r2[13]&pow|r1[9]&r2[15]&pow|r1[10]&r2[1]&sub|r1[10]&r2[15]&add|r1[11]&r2[2]&sub|r1[11]&r2[2]&pow|r1[11]&r2[6]&pow|r1[11]&r2[10]&pow|r1[11]&r2[11]&div|r1[11]&r2[14]&add|r1[11]&r2[14]&pow|r1[12]&r2[3]&sub|r1[12]&r2[13]&add|r1[13]&r2[2]&pow|r1[13]&r2[4]&sub|r1[13]&r2[6]&pow|r1[13]&r2[10]&pow|r1[13]&r2[12]&add|r1[13]&r2[13]&div|r1[13]&r2[14]&pow|r1[14]&r2[5]&sub|r1[14]&r2[11]&add|r1[15]&r2[6]&sub|r1[15]&r2[7]&div|r1[15]&r2[10]&add,
r1[0]&r2[8]&add|r1[1]&r2[7]&add|r1[1]&r2[8]&div|r1[2]&r2[3]&pow|r1[2]&r2[4]&div|r1[2]&r2[6]&add|r1[2]&r2[12]&div|r1[3]&r2[5]&add|r1[3]&r2[8]&div|r1[4]&r2[2]&div|r1[4]&r2[4]&add|r1[4]&r2[6]&div|r1[4]&r2[10]&div|r1[4]&r2[14]&div|r1[5]&r2[3]&add|r1[5]&r2[8]&div|r1[6]&r2[2]&add|r1[6]&r2[3]&pow|r1[6]&r2[4]&div|r1[6]&r2[12]&div|r1[7]&r2[1]&add|r1[7]&r2[8]&div|r1[8]&r2[0]&add|r1[8]&r2[0]&sub|r1[8]&r2[0]&mul|r1[8]&r2[1]&div|r1[8]&r2[1]&pow|r1[8]&r2[3]&div|r1[8]&r2[5]&div|r1[8]&r2[7]&div|r1[8]&r2[9]&div|r1[8]&r2[11]&div|r1[8]&r2[13]&div|r1[8]&r2[15]&div|r1[9]&r2[1]&sub|r1[9]&r2[8]&div|r1[9]&r2[15]&add|r1[10]&r2[2]&sub|r1[10]&r2[3]&pow|r1[10]&r2[4]&div|r1[10]&r2[12]&div|r1[10]&r2[14]&add|r1[11]&r2[3]&sub|r1[11]&r2[8]&div|r1[11]&r2[13]&add|r1[12]&r2[2]&div|r1[12]&r2[4]&sub|r1[12]&r2[6]&div|r1[12]&r2[10]&div|r1[12]&r2[12]&add|r1[12]&r2[14]&div|r1[13]&r2[5]&sub|r1[13]&r2[8]&div|r1[13]&r2[11]&add|r1[13]&r2[15]&pow|r1[14]&r2[3]&pow|r1[14]&r2[4]&div|r1[14]&r2[6]&sub|r1[14]&r2[10]&add|r1[14]&r2[12]&div|r1[15]&r2[7]&sub|r1[15]&r2[8]&div|r1[15]&r2[9]&add,
r1[0]&r2[7]&add|r1[1]&r2[6]&add|r1[1]&r2[7]&div|r1[2]&r2[5]&add|r1[3]&r2[4]&add|r1[3]&r2[13]&div|r1[4]&r2[3]&add|r1[5]&r2[2]&add|r1[5]&r2[11]&div|r1[6]&r2[1]&add|r1[7]&r2[0]&add|r1[7]&r2[0]&sub|r1[7]&r2[0]&mul|r1[7]&r2[1]&div|r1[7]&r2[1]&pow|r1[7]&r2[3]&pow|r1[7]&r2[5]&pow|r1[7]&r2[7]&pow|r1[7]&r2[9]&pow|r1[7]&r2[11]&pow|r1[7]&r2[13]&pow|r1[7]&r2[15]&pow|r1[8]&r2[1]&sub|r1[8]&r2[15]&add|r1[9]&r2[2]&sub|r1[9]&r2[14]&add|r1[9]&r2[15]&div|r1[10]&r2[3]&sub|r1[10]&r2[13]&add|r1[11]&r2[4]&sub|r1[11]&r2[5]&div|r1[11]&r2[12]&add|r1[12]&r2[5]&sub|r1[12]&r2[11]&add|r1[13]&r2[3]&div|r1[13]&r2[6]&sub|r1[13]&r2[10]&add|r1[14]&r2[1]&mul|r1[14]&r2[7]&sub|r1[14]&r2[9]&add|r1[15]&r2[1]&mul|r1[15]&r2[8]&add|r1[15]&r2[8]&sub|r1[15]&r2[9]&div,
r1[0]&r2[6]&add|r1[1]&r2[5]&add|r1[1]&r2[6]&div|r1[2]&r2[3]&div|r1[2]&r2[4]&add|r1[2]&r2[11]&div|r1[3]&r2[2]&div|r1[3]&r2[3]&add|r1[4]&r2[2]&add|r1[5]&r2[1]&add|r1[5]&r2[14]&div|r1[6]&r2[0]&add|r1[6]&r2[0]&sub|r1[6]&r2[0]&mul|r1[6]&r2[1]&div|r1[6]&r2[1]&pow|r1[6]&r2[9]&div|r1[7]&r2[1]&sub|r1[7]&r2[10]&div|r1[7]&r2[15]&add|r1[8]&r2[2]&sub|r1[8]&r2[14]&add|r1[9]&r2[3]&sub|r1[9]&r2[6]&div|r1[9]&r2[13]&add|r1[10]&r2[4]&sub|r1[10]&r2[7]&div|r1[10]&r2[12]&add|r1[10]&r2[15]&div|r1[11]&r2[2]&div|r1[11]&r2[5]&sub|r1[11]&r2[11]&add|r1[12]&r2[1]&mul|r1[12]&r2[6]&sub|r1[12]&r2[10]&add|r1[13]&r2[1]&mul|r1[13]&r2[7]&sub|r1[13]&r2[9]&add|r1[13]&r2[14]&div|r1[14]&r2[5]&div|r1[14]&r2[8]&add|r1[14]&r2[8]&sub|r1[14]&r2[13]&div|r1[15]&r2[7]&add|r1[15]&r2[9]&sub|r1[15]&r2[10]&div,
r1[0]&r2[5]&add|r1[1]&r2[4]&add|r1[1]&r2[5]&div|r1[2]&r2[3]&add|r1[3]&r2[2]&add|r1[3]&r2[7]&div|r1[4]&r2[1]&add|r1[5]&r2[0]&add|r1[5]&r2[0]&sub|r1[5]&r2[0]&mul|r1[5]&r2[1]&div|r1[5]&r2[1]&pow|r1[5]&r2[5]&pow|r1[5]&r2[9]&pow|r1[5]&r2[13]&pow|r1[6]&r2[1]&sub|r1[6]&r2[15]&add|r1[7]&r2[2]&sub|r1[7]&r2[3]&div|r1[7]&r2[14]&add|r1[8]&r2[3]&sub|r1[8]&r2[13]&add|r1[9]&r2[4]&sub|r1[9]&r2[12]&add|r1[9]&r2[13]&div|r1[10]&r2[1]&mul|r1[10]&r2[5]&sub|r1[10]&r2[11]&add|r1[11]&r2[1]&mul|r1[11]&r2[6]&sub|r1[11]&r2[10]&add|r1[11]&r2[15]&div|r1[12]&r2[7]&sub|r1[12]&r2[9]&add|r1[13]&r2[3]&pow|r1[13]&r2[7]&pow|r1[13]&r2[8]&add|r1[13]&r2[8]&sub|r1[13]&r2[9]&div|r1[13]&r2[11]&pow|r1[14]&r2[7]&add|r1[14]&r2[9]&sub|r1[15]&r2[2]&mul|r1[15]&r2[6]&add|r1[15]&r2[10]&sub|r1[15]&r2[11]&div,
r1[0]&r2[4]&add|r1[1]&r2[3]&add|r1[1]&r2[4]&div|r1[2]&r2[2]&add|r1[2]&r2[2]&div|r1[2]&r2[2]&pow|r1[2]&r2[10]&div|r1[3]&r2[1]&add|r1[3]&r2[12]&div|r1[4]&r2[0]&add|r1[4]&r2[0]&sub|r1[4]&r2[0]&mul|r1[4]&r2[1]&div|r1[4]&r2[1]&pow|r1[4]&r2[5]&div|r1[4]&r2[9]&div|r1[4]&r2[13]&div|r1[5]&r2[1]&sub|r1[5]&r2[4]&div|r1[5]&r2[15]&add|r1[6]&r2[2]&sub|r1[6]&r2[2]&pow|r1[6]&r2[6]&div|r1[6]&r2[14]&add|r1[6]&r2[14]&div|r1[7]&r2[3]&sub|r1[7]&r2[12]&div|r1[7]&r2[13]&add|r1[8]&r2[1]&mul|r1[8]&r2[4]&sub|r1[8]&r2[12]&add|r1[9]&r2[1]&mul|r1[9]&r2[4]&div|r1[9]&r2[5]&sub|r1[9]&r2[11]&add|r1[10]&r2[2]&div|r1[10]&r2[2]&pow|r1[10]&r2[6]&sub|r1[10]&r2[10]&add|r1[10]&r2[10]&div|r1[11]&r2[7]&sub|r1[11]&r2[9]&add|r1[11]&r2[12]&div|r1[12]&r2[2]&mul|r1[12]&r2[3]&div|r1[12]&r2[7]&div|r1[12]&r2[8]&add|r1[12]&r2[8]&sub|r1[12]&r2[11]&div|r1[12]&r2[15]&div|r1[13]&r2[2]&mul|r1[13]&r2[4]&div|r1[13]&r2[7]&add|r1[13]&r2[9]&sub|r1[14]&r2[2]&mul|r1[14]&r2[2]&pow|r1[14]&r2[6]&add|r1[14]&r2[6]&div|r1[14]&r2[10]&sub|r1[14]&r2[14]&div|r1[15]&r2[5]&add|r1[15]&r2[11]&sub|r1[15]&r2[12]&div,
r1[0]&r2[3]&add|r1[1]&r2[2]&add|r1[1]&r2[3]&div|r1[2]&r2[1]&add|r1[3]&r2[0]&add|r1[3]&r2[0]&sub|r1[3]&r2[0]&mul|r1[3]&r2[1]&div|r1[3]&r2[1]&pow|r1[3]&r2[5]&pow|r1[3]&r2[9]&pow|r1[3]&r2[13]&pow|r1[4]&r2[1]&sub|r1[4]&r2[15]&add|r1[5]&r2[2]&sub|r1[5]&r2[7]&div|r1[5]&r2[14]&add|r1[6]&r2[1]&mul|r1[6]&r2[3]&sub|r1[6]&r2[13]&add|r1[7]&r2[1]&mul|r1[7]&r2[4]&sub|r1[7]&r2[5]&div|r1[7]&r2[12]&add|r1[8]&r2[5]&sub|r1[8]&r2[11]&add|r1[9]&r2[2]&mul|r1[9]&r2[6]&sub|r1[9]&r2[10]&add|r1[9]&r2[11]&div|r1[10]&r2[2]&mul|r1[10]&r2[7]&sub|r1[10]&r2[9]&add|r1[11]&r2[2]&mul|r1[11]&r2[3]&pow|r1[11]&r2[7]&pow|r1[11]&r2[8]&add|r1[11]&r2[8]&sub|r1[11]&r2[9]&div|r1[11]&r2[11]&pow|r1[11]&r2[15]&pow|r1[12]&r2[3]&mul|r1[12]&r2[7]&add|r1[12]&r2[9]&sub|r1[13]&r2[3]&mul|r1[13]&r2[6]&add|r1[13]&r2[10]&sub|r1[13]&r2[15]&div|r1[14]&r2[3]&mul|r1[14]&r2[5]&add|r1[14]&r2[11]&sub|r1[15]&r2[3]&mul|r1[15]&r2[4]&add|r1[15]&r2[4]&mul|r1[15]&r2[12]&sub|r1[15]&r2[13]&div,
r1[0]&r2[2]&add|r1[1]&r2[1]&add|r1[1]&r2[2]&div|r1[2]&r2[0]&add|r1[2]&r2[0]&sub|r1[2]&r2[0]&mul|r1[2]&r2[1]&div|r1[2]&r2[1]&pow|r1[2]&r2[9]&div|r1[3]&r2[1]&sub|r1[3]&r2[6]&div|r1[3]&r2[15]&add|r1[4]&r2[1]&mul|r1[4]&r2[2]&sub|r1[4]&r2[14]&add|r1[5]&r2[1]&mul|r1[5]&r2[3]&sub|r1[5]&r2[10]&div|r1[5]&r2[13]&add|r1[6]&r2[2]&mul|r1[6]&r2[3]&div|r1[6]&r2[4]&sub|r1[6]&r2[11]&div|r1[6]&r2[12]&add|r1[7]&r2[2]&mul|r1[7]&r2[5]&sub|r1[7]&r2[11]&add|r1[7]&r2[14]&div|r1[8]&r2[2]&mul|r1[8]&r2[3]&mul|r1[8]&r2[6]&sub|r1[8]&r2[10]&add|r1[9]&r2[2]&div|r1[9]&r2[3]&mul|r1[9]&r2[7]&sub|r1[9]&r2[9]&add|r1[10]&r2[3]&mul|r1[10]&r2[4]&mul|r1[10]&r2[5]&div|r1[10]&r2[8]&add|r1[10]&r2[8]&sub|r1[10]&r2[13]&div|r1[11]&r2[3]&mul|r1[11]&r2[4]&mul|r1[11]&r2[6]&div|r1[11]&r2[7]&add|r1[11]&r2[9]&sub|r1[12]&r2[4]&mul|r1[12]&r2[5]&mul|r1[12]&r2[6]&add|r1[12]&r2[10]&sub|r1[13]&r2[4]&mul|r1[13]&r2[5]&add|r1[13]&r2[5]&mul|r1[13]&r2[10]&div|r1[13]&r2[11]&sub|r1[14]&r2[4]&add|r1[14]&r2[4]&mul|r1[14]&r2[5]&mul|r1[14]&r2[6]&mul|r1[14]&r2[7]&div|r1[14]&r2[12]&sub|r1[14]&r2[15]&div|r1[15]&r2[3]&add|r1[15]&r2[5]&mul|r1[15]&r2[6]&mul|r1[15]&r2[13]&sub|r1[15]&r2[14]&div,
r1[0]&r2[0]&pow|r1[0]&r2[1]&add|r1[1]&r2[0]&add|r1[1]&r2[0]&sub|r1[1]&r2[0]&mul|r1[1]&r2[0]&pow|r1[1]&r2[1]&div|r1[1]&r2[1]&pow|r1[1]&r2[2]&pow|r1[1]&r2[3]&pow|r1[1]&r2[4]&pow|r1[1]&r2[5]&pow|r1[1]&r2[6]&pow|r1[1]&r2[7]&pow|r1[1]&r2[8]&pow|r1[1]&r2[9]&pow|r1[1]&r2[10]&pow|r1[1]&r2[11]&pow|r1[1]&r2[12]&pow|r1[1]&r2[13]&pow|r1[1]&r2[14]&pow|r1[1]&r2[15]&pow|r1[2]&r2[0]&pow|r1[2]&r2[1]&sub|r1[2]&r2[1]&mul|r1[2]&r2[15]&add|r1[3]&r2[0]&pow|r1[3]&r2[1]&mul|r1[3]&r2[2]&sub|r1[3]&r2[2]&mul|r1[3]&r2[4]&pow|r1[3]&r2[8]&pow|r1[3]&r2[11]&div|r1[3]&r2[12]&pow|r1[3]&r2[14]&add|r1[4]&r2[0]&pow|r1[4]&r2[2]&mul|r1[4]&r2[3]&sub|r1[4]&r2[3]&mul|r1[4]&r2[13]&add|r1[5]&r2[0]&pow|r1[5]&r2[2]&mul|r1[5]&r2[3]&mul|r1[5]&r2[4]&sub|r1[5]&r2[4]&mul|r1[5]&r2[4]&pow|r1[5]&r2[8]&pow|r1[5]&r2[12]&add|r1[5]&r2[12]&pow|r1[5]&r2[13]&div|r1[6]&r2[0]&pow|r1[6]&r2[3]&mul|r1[6]&r2[4]&mul|r1[6]&r2[5]&sub|r1[6]&r2[5]&mul|r1[6]&r2[11]&add|r1[7]&r2[0]&pow|r1[7]&r2[2]&pow|r1[7]&r2[3]&mul|r1[7]&r2[4]&mul|r1[7]&r2[4]&pow|r1[7]&r2[5]&mul|r1[7]&r2[6]&sub|r1[7]&r2[6]&mul|r1[7]&r2[6]&pow|r1[7]&r2[7]&div|r1[7]&r2[8]&pow|r1[7]&r2[10]&add|r1[7]&r2[10]&pow|r1[7]&r2[12]&pow|r1[7]&r2[14]&pow|r1[8]&r2[0]&pow|r1[8]&r2[4]&mul|r1[8]&r2[5]&mul|r1[8]&r2[6]&mul|r1[8]&r2[7]&sub|r1[8]&r2[7]&mul|r1[8]&r2[9]&add|r1[9]&r2[0]&pow|r1[9]&r2[2]&pow|r1[9]&r2[4]&mul|r1[9]&r2[4]&pow|r1[9]&r2[5]&mul|r1[9]&r2[6]&mul|r1[9]&r2[6]&pow|r1[9]&r2[7]&mul|r1[9]&r2[8]&add|r1[9]&r2[8]&sub|r1[9]&r2[8]&mul|r1[9]&r2[8]&pow|r1[9]&r2[9]&div|r1[9]&r2[10]&pow|r1[9]&r2[12]&pow|r1[9]&r2[14]&pow|r1[10]&r2[0]&pow|r1[10]&r2[5]&mul|r1[10]&r2[6]&mul|r1[10]&r2[7]&add|r1[10]&r2[7]&mul|r1[10]&r2[8]&mul|r1[10]&r2[9]&sub|r1[10]&r2[9]&mul|r1[11]&r2[0]&pow|r1[11]&r2[3]&div|r1[11]&r2[4]&pow|r1[11]&r2[5]&mul|r1[11]&r2[6]&add|r1[11]&r2[6]&mul|r1[11]&r2[7]&mul|r1[11]&r2[8]&mul|r1[11]&r2[8]&pow|r1[11]&r2[9]&mul|r1[11]&r2[10]&sub|r1[11]&r2[10]&mul|r1[11]&r2[12]&pow|r1[12]&r2[0]&pow|r1[12]&r2[5]&add|r1[12]&r2[6]&mul|r1[12]&r2[7]&mul|r1[12]&r2[8]&mul|r1[12]&r2[9]&mul|r1[12]&r2[10]&mul|r1[12]&r2[11]&sub|r1[12]&r2[11]&mul|r1[13]&r2[0]&pow|r1[13]&r2[4]&add|r1[13]&r2[4]&pow|r1[13]&r2[5]&div|r1[13]&r2[6]&mul|r1[13]&r2[7]&mul|r1[13]&r2[8]&mul|r1[13]&r2[8]&pow|r1[13]&r2[9]&mul|r1[13]&r2[10]&mul|r1[13]&r2[11]&mul|r1[13]&r2[12]&sub|r1[13]&r2[12]&mul|r1[13]&r2[12]&pow|r1[14]&r2[0]&pow|r1[14]&r2[3]&add|r1[14]&r2[7]&mul|r1[14]&r2[8]&mul|r1[14]&r2[9]&mul|r1[14]&r2[10]&mul|r1[14]&r2[11]&mul|r1[14]&r2[12]&mul|r1[14]&r2[13]&sub|r1[14]&r2[13]&mul|r1[15]&r2[0]&pow|r1[15]&r2[2]&add|r1[15]&r2[2]&pow|r1[15]&r2[4]&pow|r1[15]&r2[6]&pow|r1[15]&r2[7]&mul|r1[15]&r2[8]&mul|r1[15]&r2[8]&pow|r1[15]&r2[9]&mul|r1[15]&r2[10]&mul|r1[15]&r2[10]&pow|r1[15]&r2[11]&mul|r1[15]&r2[12]&mul|r1[15]&r2[12]&pow|r1[15]&r2[13]&mul|r1[15]&r2[14]&sub|r1[15]&r2[14]&mul|r1[15]&r2[15]&div,
r1[0]&r2[0]&add|r1[0]&r2[0]&sub|r1[0]&r2[0]&div|r1[0]&r2[0]&mul|r1[0]&r2[0]&act_func|r1[0]&r2[0]&act_func_2_1|r1[0]&r2[1]&sub|r1[0]&r2[1]&div|r1[0]&r2[1]&mul|r1[0]&r2[1]&pow|r1[0]&r2[1]&act_func|r1[0]&r2[1]&act_func_2_1|r1[0]&r2[2]&sub|r1[0]&r2[2]&div|r1[0]&r2[2]&mul|r1[0]&r2[2]&pow|r1[0]&r2[2]&act_func|r1[0]&r2[2]&act_func_2_1|r1[0]&r2[3]&sub|r1[0]&r2[3]&div|r1[0]&r2[3]&mul|r1[0]&r2[3]&pow|r1[0]&r2[3]&act_func|r1[0]&r2[3]&act_func_2_1|r1[0]&r2[4]&sub|r1[0]&r2[4]&div|r1[0]&r2[4]&mul|r1[0]&r2[4]&pow|r1[0]&r2[4]&act_func|r1[0]&r2[4]&act_func_2_1|r1[0]&r2[5]&sub|r1[0]&r2[5]&div|r1[0]&r2[5]&mul|r1[0]&r2[5]&pow|r1[0]&r2[5]&act_func|r1[0]&r2[5]&act_func_2_1|r1[0]&r2[6]&sub|r1[0]&r2[6]&div|r1[0]&r2[6]&mul|r1[0]&r2[6]&pow|r1[0]&r2[6]&act_func|r1[0]&r2[6]&act_func_2_1|r1[0]&r2[7]&sub|r1[0]&r2[7]&div|r1[0]&r2[7]&mul|r1[0]&r2[7]&pow|r1[0]&r2[7]&act_func|r1[0]&r2[7]&act_func_2_1|r1[0]&r2[8]&sub|r1[0]&r2[8]&div|r1[0]&r2[8]&mul|r1[0]&r2[8]&pow|r1[0]&r2[8]&act_func|r1[0]&r2[8]&act_func_2_1|r1[0]&r2[9]&sub|r1[0]&r2[9]&div|r1[0]&r2[9]&mul|r1[0]&r2[9]&pow|r1[0]&r2[9]&act_func|r1[0]&r2[9]&act_func_2_1|r1[0]&r2[10]&sub|r1[0]&r2[10]&div|r1[0]&r2[10]&mul|r1[0]&r2[10]&pow|r1[0]&r2[10]&act_func|r1[0]&r2[10]&act_func_2_1|r1[0]&r2[11]&sub|r1[0]&r2[11]&div|r1[0]&r2[11]&mul|r1[0]&r2[11]&pow|r1[0]&r2[11]&act_func|r1[0]&r2[11]&act_func_2_1|r1[0]&r2[12]&sub|r1[0]&r2[12]&div|r1[0]&r2[12]&mul|r1[0]&r2[12]&pow|r1[0]&r2[12]&act_func|r1[0]&r2[12]&act_func_2_1|r1[0]&r2[13]&sub|r1[0]&r2[13]&div|r1[0]&r2[13]&mul|r1[0]&r2[13]&pow|r1[0]&r2[13]&act_func|r1[0]&r2[13]&act_func_2_1|r1[0]&r2[14]&sub|r1[0]&r2[14]&div|r1[0]&r2[14]&mul|r1[0]&r2[14]&pow|r1[0]&r2[14]&act_func|r1[0]&r2[14]&act_func_2_1|r1[0]&r2[15]&sub|r1[0]&r2[15]&div|r1[0]&r2[15]&mul|r1[0]&r2[15]&pow|r1[0]&r2[15]&act_func|r1[0]&r2[15]&act_func_2_1|r1[1]&r2[0]&div|r1[1]&r2[0]&act_func|r1[1]&r2[0]&act_func_2_1|r1[1]&r2[1]&sub|r1[1]&r2[1]&mul|r1[1]&r2[1]&act_func|r1[1]&r2[1]&act_func_2_1|r1[1]&r2[2]&sub|r1[1]&r2[2]&mul|r1[1]&r2[2]&act_func|r1[1]&r2[2]&act_func_2_1|r1[1]&r2[3]&sub|r1[1]&r2[3]&mul|r1[1]&r2[3]&act_func|r1[1]&r2[3]&act_func_2_1|r1[1]&r2[4]&sub|r1[1]&r2[4]&mul|r1[1]&r2[4]&act_func|r1[1]&r2[4]&act_func_2_1|r1[1]&r2[5]&sub|r1[1]&r2[5]&mul|r1[1]&r2[5]&act_func|r1[1]&r2[5]&act_func_2_1|r1[1]&r2[6]&sub|r1[1]&r2[6]&mul|r1[1]&r2[6]&act_func|r1[1]&r2[6]&act_func_2_1|r1[1]&r2[7]&sub|r1[1]&r2[7]&mul|r1[1]&r2[7]&act_func|r1[1]&r2[7]&act_func_2_1|r1[1]&r2[8]&sub|r1[1]&r2[8]&mul|r1[1]&r2[8]&act_func|r1[1]&r2[8]&act_func_2_1|r1[1]&r2[9]&sub|r1[1]&r2[9]&mul|r1[1]&r2[9]&act_func|r1[1]&r2[9]&act_func_2_1|r1[1]&r2[10]&sub|r1[1]&r2[10]&mul|r1[1]&r2[10]&act_func|r1[1]&r2[10]&act_func_2_1|r1[1]&r2[11]&sub|r1[1]&r2[11]&mul|r1[1]&r2[11]&act_func|r1[1]&r2[11]&act_func_2_1|r1[1]&r2[12]&sub|r1[1]&r2[12]&mul|r1[1]&r2[12]&act_func|r1[1]&r2[12]&act_func_2_1|r1[1]&r2[13]&sub|r1[1]&r2[13]&mul|r1[1]&r2[13]&act_func|r1[1]&r2[13]&act_func_2_1|r1[1]&r2[14]&sub|r1[1]&r2[14]&mul|r1[1]&r2[14]&act_func|r1[1]&r2[14]&act_func_2_1|r1[1]&r2[15]&add|r1[1]&r2[15]&sub|r1[1]&r2[15]&mul|r1[1]&r2[15]&act_func|r1[1]&r2[15]&act_func_2_1|r1[2]&r2[0]&div|r1[2]&r2[0]&act_func|r1[2]&r2[0]&act_func_2_1|r1[2]&r2[1]&act_func|r1[2]&r2[1]&act_func_2_1|r1[2]&r2[2]&sub|r1[2]&r2[2]&mul|r1[2]&r2[2]&act_func|r1[2]&r2[2]&act_func_2_1|r1[2]&r2[3]&sub|r1[2]&r2[3]&mul|r1[2]&r2[3]&act_func|r1[2]&r2[3]&act_func_2_1|r1[2]&r2[4]&sub|r1[2]&r2[4]&mul|r1[2]&r2[4]&pow|r1[2]&r2[4]&act_func|r1[2]&r2[4]&act_func_2_1|r1[2]&r2[5]&sub|r1[2]&r2[5]&mul|r1[2]&r2[5]&pow|r1[2]&r2[5]&act_func|r1[2]&r2[5]&act_func_2_1|r1[2]&r2[6]&sub|r1[2]&r2[6]&mul|r1[2]&r2[6]&pow|r1[2]&r2[6]&act_func|r1[2]&r2[6]&act_func_2_1|r1[2]&r2[7]&sub|r1[2]&r2[7]&mul|r1[2]&r2[7]&pow|r1[2]&r2[7]&act_func|r1[2]&r2[7]&act_func_2_1|r1[2]&r2[8]&sub|r1[2]&r2[8]&div|r1[2]&r2[8]&mul|r1[2]&r2[8]&pow|r1[2]&r2[8]&act_func|r1[2]&r2[8]&act_func_2_1|r1[2]&r2[9]&sub|r1[2]&r2[9]&mul|r1[2]&r2[9]&pow|r1[2]&r2[9]&act_func|r1[2]&r2[9]&act_func_2_1|r1[2]&r2[10]&sub|r1[2]&r2[10]&mul|r1[2]&r2[10]&pow|r1[2]&r2[10]&act_func|r1[2]&r2[10]&act_func_2_1|r1[2]&r2[11]&sub|r1[2]&r2[11]&mul|r1[2]&r2[11]&pow|r1[2]&r2[11]&act_func|r1[2]&r2[11]&act_func_2_1|r1[2]&r2[12]&sub|r1[2]&r2[12]&mul|r1[2]&r2[12]&pow|r1[2]&r2[12]&act_func|r1[2]&r2[12]&act_func_2_1|r1[2]&r2[13]&sub|r1[2]&r2[13]&mul|r1[2]&r2[13]&pow|r1[2]&r2[13]&act_func|r1[2]&r2[13]&act_func_2_1|r1[2]&r2[14]&add|r1[2]&r2[14]&sub|r1[2]&r2[14]&mul|r1[2]&r2[14]&pow|r1[2]&r2[14]&act_func|r1[2]&r2[14]&act_func_2_1|r1[2]&r2[15]&sub|r1[2]&r2[15]&mul|r1[2]&r2[15]&pow|r1[2]&r2[15]&act_func|r1[2]&r2[15]&act_func_2_1|r1[3]&r2[0]&div|r1[3]&r2[0]&act_func|r1[3]&r2[0]&act_func_2_1|r1[3]&r2[1]&act_func|r1[3]&r2[1]&act_func_2_1|r1[3]&r2[2]&act_func|r1[3]&r2[2]&act_func_2_1|r1[3]&r2[3]&sub|r1[3]&r2[3]&mul|r1[3]&r2[3]&act_func|r1[3]&r2[3]&act_func_2_1|r1[3]&r2[4]&sub|r1[3]&r2[4]&mul|r1[3]&r2[4]&act_func|r1[3]&r2[4]&act_func_2_1|r1[3]&r2[5]&sub|r1[3]&r2[5]&mul|r1[3]&r2[5]&act_func|r1[3]&r2[5]&act_func_2_1|r1[3]&r2[6]&sub|r1[3]&r2[6]&mul|r1[3]&r2[6]&act_func|r1[3]&r2[6]&act_func_2_1|r1[3]&r2[7]&sub|r1[3]&r2[7]&mul|r1[3]&r2[7]&act_func|r1[3]&r2[7]&act_func_2_1|r1[3]&r2[8]&sub|r1[3]&r2[8]&mul|r1[3]&r2[8]&act_func|r1[3]&r2[8]&act_func_2_1|r1[3]&r2[9]&sub|r1[3]&r2[9]&mul|r1[3]&r2[9]&act_func|r1[3]&r2[9]&act_func_2_1|r1[3]&r2[10]&sub|r1[3]&r2[10]&mul|r1[3]&r2[10]&act_func|r1[3]&r2[10]&act_func_2_1|r1[3]&r2[11]&sub|r1[3]&r2[11]&mul|r1[3]&r2[11]&act_func|r1[3]&r2[11]&act_func_2_1|r1[3]&r2[12]&sub|r1[3]&r2[12]&mul|r1[3]&r2[12]&act_func|r1[3]&r2[12]&act_func_2_1|r1[3]&r2[13]&add|r1[3]&r2[13]&sub|r1[3]&r2[13]&mul|r1[3]&r2[13]&act_func|r1[3]&r2[13]&act_func_2_1|r1[3]&r2[14]&sub|r1[3]&r2[14]&mul|r1[3]&r2[14]&act_func|r1[3]&r2[14]&act_func_2_1|r1[3]&r2[15]&sub|r1[3]&r2[15]&mul|r1[3]&r2[15]&act_func|r1[3]&r2[15]&act_func_2_1|r1[4]&r2[0]&div|r1[4]&r2[0]&act_func|r1[4]&r2[0]&act_func_2_1|r1[4]&r2[1]&act_func|r1[4]&r2[1]&act_func_2_1|r1[4]&r2[2]&pow|r1[4]&r2[2]&act_func|r1[4]&r2[2]&act_func_2_1|r1[4]&r2[3]&pow|r1[4]&r2[3]&act_func|r1[4]&r2[3]&act_func_2_1|r1[4]&r2[4]&sub|r1[4]&r2[4]&div|r1[4]&r2[4]&mul|r1[4]&r2[4]&pow|r1[4]&r2[4]&act_func|r1[4]&r2[4]&act_func_2_1|r1[4]&r2[5]&sub|r1[4]&r2[5]&mul|r1[4]&r2[5]&pow|r1[4]&r2[5]&act_func|r1[4]&r2[5]&act_func_2_1|r1[4]&r2[6]&sub|r1[4]&r2[6]&mul|r1[4]&r2[6]&pow|r1[4]&r2[6]&act_func|r1[4]&r2[6]&act_func_2_1|r1[4]&r2[7]&sub|r1[4]&r2[7]&mul|r1[4]&r2[7]&pow|r1[4]&r2[7]&act_func|r1[4]&r2[7]&act_func_2_1|r1[4]&r2[8]&sub|r1[4]&r2[8]&div|r1[4]&r2[8]&mul|r1[4]&r2[8]&pow|r1[4]&r2[8]&act_func|r1[4]&r2[8]&act_func_2_1|r1[4]&r2[9]&sub|r1[4]&r2[9]&mul|r1[4]&r2[9]&pow|r1[4]&r2[9]&act_func|r1[4]&r2[9]&act_func_2_1|r1[4]&r2[10]&sub|r1[4]&r2[10]&mul|r1[4]&r2[10]&pow|r1[4]&r2[10]&act_func|r1[4]&r2[10]&act_func_2_1|r1[4]&r2[11]&sub|r1[4]&r2[11]&mul|r1[4]&r2[11]&pow|r1[4]&r2[11]&act_func|r1[4]&r2[11]&act_func_2_1|r1[4]&r2[12]&add|r1[4]&r2[12]&sub|r1[4]&r2[12]&div|r1[4]&r2[12]&mul|r1[4]&r2[12]&pow|r1[4]&r2[12]&act_func|r1[4]&r2[12]&act_func_2_1|r1[4]&r2[13]&sub|r1[4]&r2[13]&mul|r1[4]&r2[13]&pow|r1[4]&r2[13]&act_func|r1[4]&r2[13]&act_func_2_1|r1[4]&r2[14]&sub|r1[4]&r2[14]&mul|r1[4]&r2[14]&pow|r1[4]&r2[14]&act_func|r1[4]&r2[14]&act_func_2_1|r1[4]&r2[15]&sub|r1[4]&r2[15]&mul|r1[4]&r2[15]&pow|r1[4]&r2[15]&act_func|r1[4]&r2[15]&act_func_2_1|r1[5]&r2[0]&div|r1[5]&r2[0]&act_func|r1[5]&r2[0]&act_func_2_1|r1[5]&r2[1]&act_func|r1[5]&r2[1]&act_func_2_1|r1[5]&r2[2]&act_func|r1[5]&r2[2]&act_func_2_1|r1[5]&r2[3]&act_func|r1[5]&r2[3]&act_func_2_1|r1[5]&r2[4]&act_func|r1[5]&r2[4]&act_func_2_1|r1[5]&r2[5]&sub|r1[5]&r2[5]&mul|r1[5]&r2[5]&act_func|r1[5]&r2[5]&act_func_2_1|r1[5]&r2[6]&sub|r1[5]&r2[6]&mul|r1[5]&r2[6]&act_func|r1[5]&r2[6]&act_func_2_1|r1[5]&r2[7]&sub|r1[5]&r2[7]&mul|r1[5]&r2[7]&act_func|r1[5]&r2[7]&act_func_2_1|r1[5]&r2[8]&sub|r1[5]&r2[8]&mul|r1[5]&r2[8]&act_func|r1[5]&r2[8]&act_func_2_1|r1[5]&r2[9]&sub|r1[5]&r2[9]&mul|r1[5]&r2[9]&act_func|r1[5]&r2[9]&act_func_2_1|r1[5]&r2[10]&sub|r1[5]&r2[10]&mul|r1[5]&r2[10]&act_func|r1[5]&r2[10]&act_func_2_1|r1[5]&r2[11]&add|r1[5]&r2[11]&sub|r1[5]&r2[11]&mul|r1[5]&r2[11]&act_func|r1[5]&r2[11]&act_func_2_1|r1[5]&r2[12]&sub|r1[5]&r2[12]&mul|r1[5]&r2[12]&act_func|r1[5]&r2[12]&act_func_2_1|r1[5]&r2[13]&sub|r1[5]&r2[13]&mul|r1[5]&r2[13]&act_func|r1[5]&r2[13]&act_func_2_1|r1[5]&r2[14]&sub|r1[5]&r2[14]&mul|r1[5]&r2[14]&act_func|r1[5]&r2[14]&act_func_2_1|r1[5]&r2[15]&sub|r1[5]&r2[15]&mul|r1[5]&r2[15]&act_func|r1[5]&r2[15]&act_func_2_1|r1[6]&r2[0]&div|r1[6]&r2[0]&act_func|r1[6]&r2[0]&act_func_2_1|r1[6]&r2[1]&act_func|r1[6]&r2[1]&act_func_2_1|r1[6]&r2[2]&act_func|r1[6]&r2[2]&act_func_2_1|r1[6]&r2[3]&act_func|r1[6]&r2[3]&act_func_2_1|r1[6]&r2[4]&pow|r1[6]&r2[4]&act_func|r1[6]&r2[4]&act_func_2_1|r1[6]&r2[5]&pow|r1[6]&r2[5]&act_func|r1[6]&r2[5]&act_func_2_1|r1[6]&r2[6]&sub|r1[6]&r2[6]&mul|r1[6]&r2[6]&pow|r1[6]&r2[6]&act_func|r1[6]&r2[6]&act_func_2_1|r1[6]&r2[7]&sub|r1[6]&r2[7]&mul|r1[6]&r2[7]&pow|r1[6]&r2[7]&act_func|r1[6]&r2[7]&act_func_2_1|r1[6]&r2[8]&sub|r1[6]&r2[8]&div|r1[6]&r2[8]&mul|r1[6]&r2[8]&pow|r1[6]&r2[8]&act_func|r1[6]&r2[8]&act_func_2_1|r1[6]&r2[9]&sub|r1[6]&r2[9]&mul|r1[6]&r2[9]&pow|r1[6]&r2[9]&act_func|r1[6]&r2[9]&act_func_2_1|r1[6]&r2[10]&add|r1[6]&r2[10]&sub|r1[6]&r2[10]&mul|r1[6]&r2[10]&pow|r1[6]&r2[10]&act_func|r1[6]&r2[10]&act_func_2_1|r1[6]&r2[11]&sub|r1[6]&r2[11]&mul|r1[6]&r2[11]&pow|r1[6]&r2[11]&act_func|r1[6]&r2[11]&act_func_2_1|r1[6]&r2[12]&sub|r1[6]&r2[12]&mul|r1[6]&r2[12]&pow|r1[6]&r2[12]&act_func|r1[6]&r2[12]&act_func_2_1|r1[6]&r2[13]&sub|r1[6]&r2[13]&mul|r1[6]&r2[13]&pow|r1[6]&r2[13]&act_func|r1[6]&r2[13]&act_func_2_1|r1[6]&r2[14]&sub|r1[6]&r2[14]&mul|r1[6]&r2[14]&pow|r1[6]&r2[14]&act_func|r1[6]&r2[14]&act_func_2_1|r1[6]&r2[15]&sub|r1[6]&r2[15]&mul|r1[6]&r2[15]&pow|r1[6]&r2[15]&act_func|r1[6]&r2[15]&act_func_2_1|r1[7]&r2[0]&div|r1[7]&r2[0]&act_func|r1[7]&r2[0]&act_func_2_1|r1[7]&r2[1]&act_func|r1[7]&r2[1]&act_func_2_1|r1[7]&r2[2]&act_func|r1[7]&r2[2]&act_func_2_1|r1[7]&r2[3]&act_func|r1[7]&r2[3]&act_func_2_1|r1[7]&r2[4]&act_func|r1[7]&r2[4]&act_func_2_1|r1[7]&r2[5]&act_func|r1[7]&r2[5]&act_func_2_1|r1[7]&r2[6]&act_func|r1[7]&r2[6]&act_func_2_1|r1[7]&r2[7]&sub|r1[7]&r2[7]&mul|r1[7]&r2[7]&act_func|r1[7]&r2[7]&act_func_2_1|r1[7]&r2[8]&sub|r1[7]&r2[8]&mul|r1[7]&r2[8]&act_func|r1[7]&r2[8]&act_func_2_1|r1[7]&r2[9]&add|r1[7]&r2[9]&sub|r1[7]&r2[9]&mul|r1[7]&r2[9]&act_func|r1[7]&r2[9]&act_func_2_1|r1[7]&r2[10]&sub|r1[7]&r2[10]&mul|r1[7]&r2[10]&act_func|r1[7]&r2[10]&act_func_2_1|r1[7]&r2[11]&sub|r1[7]&r2[11]&mul|r1[7]&r2[11]&act_func|r1[7]&r2[11]&act_func_2_1|r1[7]&r2[12]&sub|r1[7]&r2[12]&mul|r1[7]&r2[12]&act_func|r1[7]&r2[12]&act_func_2_1|r1[7]&r2[13]&sub|r1[7]&r2[13]&mul|r1[7]&r2[13]&act_func|r1[7]&r2[13]&act_func_2_1|r1[7]&r2[14]&sub|r1[7]&r2[14]&mul|r1[7]&r2[14]&act_func|r1[7]&r2[14]&act_func_2_1|r1[7]&r2[15]&sub|r1[7]&r2[15]&mul|r1[7]&r2[15]&act_func|r1[7]&r2[15]&act_func_2_1|r1[8]&r2[0]&div|r1[8]&r2[0]&act_func|r1[8]&r2[0]&act_func_2_1|r1[8]&r2[1]&act_func|r1[8]&r2[1]&act_func_2_1|r1[8]&r2[2]&div|r1[8]&r2[2]&pow|r1[8]&r2[2]&act_func|r1[8]&r2[2]&act_func_2_1|r1[8]&r2[3]&pow|r1[8]&r2[3]&act_func|r1[8]&r2[3]&act_func_2_1|r1[8]&r2[4]&div|r1[8]&r2[4]&pow|r1[8]&r2[4]&act_func|r1[8]&r2[4]&act_func_2_1|r1[8]&r2[5]&pow|r1[8]&r2[5]&act_func|r1[8]&r2[5]&act_func_2_1|r1[8]&r2[6]&div|r1[8]&r2[6]&pow|r1[8]&r2[6]&act_func|r1[8]&r2[6]&act_func_2_1|r1[8]&r2[7]&pow|r1[8]&r2[7]&act_func|r1[8]&r2[7]&act_func_2_1|r1[8]&r2[8]&add|r1[8]&r2[8]&sub|r1[8]&r2[8]&div|r1[8]&r2[8]&mul|r1[8]&r2[8]&pow|r1[8]&r2[8]&act_func|r1[8]&r2[8]&act_func_2_1|r1[8]&r2[9]&sub|r1[8]&r2[9]&mul|r1[8]&r2[9]&pow|r1[8]&r2[9]&act_func|r1[8]&r2[9]&act_func_2_1|r1[8]&r2[10]&sub|r1[8]&r2[10]&div|r1[8]&r2[10]&mul|r1[8]&r2[10]&pow|r1[8]&r2[10]&act_func|r1[8]&r2[10]&act_func_2_1|r1[8]&r2[11]&sub|r1[8]&r2[11]&mul|r1[8]&r2[11]&pow|r1[8]&r2[11]&act_func|r1[8]&r2[11]&act_func_2_1|r1[8]&r2[12]&sub|r1[8]&r2[12]&div|r1[8]&r2[12]&mul|r1[8]&r2[12]&pow|r1[8]&r2[12]&act_func|r1[8]&r2[12]&act_func_2_1|r1[8]&r2[13]&sub|r1[8]&r2[13]&mul|r1[8]&r2[13]&pow|r1[8]&r2[13]&act_func|r1[8]&r2[13]&act_func_2_1|r1[8]&r2[14]&sub|r1[8]&r2[14]&div|r1[8]&r2[14]&mul|r1[8]&r2[14]&pow|r1[8]&r2[14]&act_func|r1[8]&r2[14]&act_func_2_1|r1[8]&r2[15]&sub|r1[8]&r2[15]&mul|r1[8]&r2[15]&pow|r1[8]&r2[15]&act_func|r1[8]&r2[15]&act_func_2_1|r1[9]&r2[0]&div|r1[9]&r2[0]&act_func|r1[9]&r2[0]&act_func_2_1|r1[9]&r2[1]&act_func|r1[9]&r2[1]&act_func_2_1|r1[9]&r2[2]&act_func|r1[9]&r2[2]&act_func_2_1|r1[9]&r2[3]&act_func|r1[9]&r2[3]&act_func_2_1|r1[9]&r2[4]&act_func|r1[9]&r2[4]&act_func_2_1|r1[9]&r2[5]&act_func|r1[9]&r2[5]&act_func_2_1|r1[9]&r2[6]&act_func|r1[9]&r2[6]&act_func_2_1|r1[9]&r2[7]&add|r1[9]&r2[7]&act_func|r1[9]&r2[7]&act_func_2_1|r1[9]&r2[8]&act_func|r1[9]&r2[8]&act_func_2_1|r1[9]&r2[9]&sub|r1[9]&r2[9]&mul|r1[9]&r2[9]&act_func|r1[9]&r2[9]&act_func_2_1|r1[9]&r2[10]&sub|r1[9]&r2[10]&mul|r1[9]&r2[10]&act_func|r1[9]&r2[10]&act_func_2_1|r1[9]&r2[11]&sub|r1[9]&r2[11]&mul|r1[9]&r2[11]&act_func|r1[9]&r2[11]&act_func_2_1|r1[9]&r2[12]&sub|r1[9]&r2[12]&mul|r1[9]&r2[12]&act_func|r1[9]&r2[12]&act_func_2_1|r1[9]&r2[13]&sub|r1[9]&r2[13]&mul|r1[9]&r2[13]&act_func|r1[9]&r2[13]&act_func_2_1|r1[9]&r2[14]&sub|r1[9]&r2[14]&mul|r1[9]&r2[14]&act_func|r1[9]&r2[14]&act_func_2_1|r1[9]&r2[15]&sub|r1[9]&r2[15]&mul|r1[9]&r2[15]&act_func|r1[9]&r2[15]&act_func_2_1|r1[10]&r2[0]&div|r1[10]&r2[0]&act_func|r1[10]&r2[0]&act_func_2_1|r1[10]&r2[1]&act_func|r1[10]&r2[1]&act_func_2_1|r1[10]&r2[2]&act_func|r1[10]&r2[2]&act_func_2_1|r1[10]&r2[3]&act_func|r1[10]&r2[3]&act_func_2_1|r1[10]&r2[4]&pow|r1[10]&r2[4]&act_func|r1[10]&r2[4]&act_func_2_1|r1[10]&r2[5]&pow|r1[10]&r2[5]&act_func|r1[10]&r2[5]&act_func_2_1|r1[10]&r2[6]&add|r1[10]&r2[6]&pow|r1[10]&r2[6]&act_func|r1[10]&r2[6]&act_func_2_1|r1[10]&r2[7]&pow|r1[10]&r2[7]&act_func|r1[10]&r2[7]&act_func_2_1|r1[10]&r2[8]&div|r1[10]&r2[8]&pow|r1[10]&r2[8]&act_func|r1[10]&r2[8]&act_func_2_1|r1[10]&r2[9]&pow|r1[10]&r2[9]&act_func|r1[10]&r2[9]&act_func_2_1|r1[10]&r2[10]&sub|r1[10]&r2[10]&mul|r1[10]&r2[10]&pow|r1[10]&r2[10]&act_func|r1[10]&r2[10]&act_func_2_1|r1[10]&r2[11]&sub|r1[10]&r2[11]&mul|r1[10]&r2[11]&pow|r1[10]&r2[11]&act_func|r1[10]&r2[11]&act_func_2_1|r1[10]&r2[12]&sub|r1[10]&r2[12]&mul|r1[10]&r2[12]&pow|r1[10]&r2[12]&act_func|r1[10]&r2[12]&act_func_2_1|r1[10]&r2[13]&sub|r1[10]&r2[13]&mul|r1[10]&r2[13]&pow|r1[10]&r2[13]&act_func|r1[10]&r2[13]&act_func_2_1|r1[10]&r2[14]&sub|r1[10]&r2[14]&mul|r1[10]&r2[14]&pow|r1[10]&r2[14]&act_func|r1[10]&r2[14]&act_func_2_1|r1[10]&r2[15]&sub|r1[10]&r2[15]&mul|r1[10]&r2[15]&pow|r1[10]&r2[15]&act_func|r1[10]&r2[15]&act_func_2_1|r1[11]&r2[0]&div|r1[11]&r2[0]&act_func|r1[11]&r2[0]&act_func_2_1|r1[11]&r2[1]&act_func|r1[11]&r2[1]&act_func_2_1|r1[11]&r2[2]&act_func|r1[11]&r2[2]&act_func_2_1|r1[11]&r2[3]&act_func|r1[11]&r2[3]&act_func_2_1|r1[11]&r2[4]&act_func|r1[11]&r2[4]&act_func_2_1|r1[11]&r2[5]&add|r1[11]&r2[5]&act_func|r1[11]&r2[5]&act_func_2_1|r1[11]&r2[6]&act_func|r1[11]&r2[6]&act_func_2_1|r1[11]&r2[7]&act_func|r1[11]&r2[7]&act_func_2_1|r1[11]&r2[8]&act_func|r1[11]&r2[8]&act_func_2_1|r1[11]&r2[9]&act_func|r1[11]&r2[9]&act_func_2_1|r1[11]&r2[10]&act_func|r1[11]&r2[10]&act_func_2_1|r1[11]&r2[11]&sub|r1[11]&r2[11]&mul|r1[11]&r2[11]&act_func|r1[11]&r2[11]&act_func_2_1|r1[11]&r2[12]&sub|r1[11]&r2[12]&mul|r1[11]&r2[12]&act_func|r1[11]&r2[12]&act_func_2_1|r1[11]&r2[13]&sub|r1[11]&r2[13]&mul|r1[11]&r2[13]&act_func|r1[11]&r2[13]&act_func_2_1|r1[11]&r2[14]&sub|r1[11]&r2[14]&mul|r1[11]&r2[14]&act_func|r1[11]&r2[14]&act_func_2_1|r1[11]&r2[15]&sub|r1[11]&r2[15]&mul|r1[11]&r2[15]&act_func|r1[11]&r2[15]&act_func_2_1|r1[12]&r2[0]&div|r1[12]&r2[0]&act_func|r1[12]&r2[0]&act_func_2_1|r1[12]&r2[1]&act_func|r1[12]&r2[1]&act_func_2_1|r1[12]&r2[2]&pow|r1[12]&r2[2]&act_func|r1[12]&r2[2]&act_func_2_1|r1[12]&r2[3]&pow|r1[12]&r2[3]&act_func|r1[12]&r2[3]&act_func_2_1|r1[12]&r2[4]&add|r1[12]&r2[4]&div|r1[12]&r2[4]&pow|r1[12]&r2[4]&act_func|r1[12]&r2[4]&act_func_2_1|r1[12]&r2[5]&pow|r1[12]&r2[5]&act_func|r1[12]&r2[5]&act_func_2_1|r1[12]&r2[6]&pow|r1[12]&r2[6]&act_func|r1[12]&r2[6]&act_func_2_1|r1[12]&r2[7]&pow|r1[12]&r2[7]&act_func|r1[12]&r2[7]&act_func_2_1|r1[12]&r2[8]&div|r1[12]&r2[8]&pow|r1[12]&r2[8]&act_func|r1[12]&r2[8]&act_func_2_1|r1[12]&r2[9]&pow|r1[12]&r2[9]&act_func|r1[12]&r2[9]&act_func_2_1|r1[12]&r2[10]&pow|r1[12]&r2[10]&act_func|r1[12]&r2[10]&act_func_2_1|r1[12]&r2[11]&pow|r1[12]&r2[11]&act_func|r1[12]&r2[11]&act_func_2_1|r1[12]&r2[12]&sub|r1[12]&r2[12]&div|r1[12]&r2[12]&mul|r1[12]&r2[12]&pow|r1[12]&r2[12]&act_func|r1[12]&r2[12]&act_func_2_1|r1[12]&r2[13]&sub|r1[12]&r2[13]&mul|r1[12]&r2[13]&pow|r1[12]&r2[13]&act_func|r1[12]&r2[13]&act_func_2_1|r1[12]&r2[14]&sub|r1[12]&r2[14]&mul|r1[12]&r2[14]&pow|r1[12]&r2[14]&act_func|r1[12]&r2[14]&act_func_2_1|r1[12]&r2[15]&sub|r1[12]&r2[15]&mul|r1[12]&r2[15]&pow|r1[12]&r2[15]&act_func|r1[12]&r2[15]&act_func_2_1|r1[13]&r2[0]&div|r1[13]&r2[0]&act_func|r1[13]&r2[0]&act_func_2_1|r1[13]&r2[1]&act_func|r1[13]&r2[1]&act_func_2_1|r1[13]&r2[2]&act_func|r1[13]&r2[2]&act_func_2_1|r1[13]&r2[3]&add|r1[13]&r2[3]&act_func|r1[13]&r2[3]&act_func_2_1|r1[13]&r2[4]&act_func|r1[13]&r2[4]&act_func_2_1|r1[13]&r2[5]&act_func|r1[13]&r2[5]&act_func_2_1|r1[13]&r2[6]&act_func|r1[13]&r2[6]&act_func_2_1|r1[13]&r2[7]&act_func|r1[13]&r2[7]&act_func_2_1|r1[13]&r2[8]&act_func|r1[13]&r2[8]&act_func_2_1|r1[13]&r2[9]&act_func|r1[13]&r2[9]&act_func_2_1|r1[13]&r2[10]&act_func|r1[13]&r2[10]&act_func_2_1|r1[13]&r2[11]&act_func|r1[13]&r2[11]&act_func_2_1|r1[13]&r2[12]&act_func|r1[13]&r2[12]&act_func_2_1|r1[13]&r2[13]&sub|r1[13]&r2[13]&mul|r1[13]&r2[13]&act_func|r1[13]&r2[13]&act_func_2_1|r1[13]&r2[14]&sub|r1[13]&r2[14]&mul|r1[13]&r2[14]&act_func|r1[13]&r2[14]&act_func_2_1|r1[13]&r2[15]&sub|r1[13]&r2[15]&mul|r1[13]&r2[15]&act_func|r1[13]&r2[15]&act_func_2_1|r1[14]&r2[0]&div|r1[14]&r2[0]&act_func|r1[14]&r2[0]&act_func_2_1|r1[14]&r2[1]&act_func|r1[14]&r2[1]&act_func_2_1|r1[14]&r2[2]&add|r1[14]&r2[2]&act_func|r1[14]&r2[2]&act_func_2_1|r1[14]&r2[3]&act_func|r1[14]&r2[3]&act_func_2_1|r1[14]&r2[4]&pow|r1[14]&r2[4]&act_func|r1[14]&r2[4]&act_func_2_1|r1[14]&r2[5]&pow|r1[14]&r2[5]&act_func|r1[14]&r2[5]&act_func_2_1|r1[14]&r2[6]&pow|r1[14]&r2[6]&act_func|r1[14]&r2[6]&act_func_2_1|r1[14]&r2[7]&pow|r1[14]&r2[7]&act_func|r1[14]&r2[7]&act_func_2_1|r1[14]&r2[8]&div|r1[14]&r2[8]&pow|r1[14]&r2[8]&act_func|r1[14]&r2[8]&act_func_2_1|r1[14]&r2[9]&pow|r1[14]&r2[9]&act_func|r1[14]&r2[9]&act_func_2_1|r1[14]&r2[10]&pow|r1[14]&r2[10]&act_func|r1[14]&r2[10]&act_func_2_1|r1[14]&r2[11]&pow|r1[14]&r2[11]&act_func|r1[14]&r2[11]&act_func_2_1|r1[14]&r2[12]&pow|r1[14]&r2[12]&act_func|r1[14]&r2[12]&act_func_2_1|r1[14]&r2[13]&pow|r1[14]&r2[13]&act_func|r1[14]&r2[13]&act_func_2_1|r1[14]&r2[14]&sub|r1[14]&r2[14]&mul|r1[14]&r2[14]&pow|r1[14]&r2[14]&act_func|r1[14]&r2[14]&act_func_2_1|r1[14]&r2[15]&sub|r1[14]&r2[15]&mul|r1[14]&r2[15]&pow|r1[14]&r2[15]&act_func|r1[14]&r2[15]&act_func_2_1|r1[15]&r2[0]&div|r1[15]&r2[0]&act_func|r1[15]&r2[0]&act_func_2_1|r1[15]&r2[1]&add|r1[15]&r2[1]&act_func|r1[15]&r2[1]&act_func_2_1|r1[15]&r2[2]&act_func|r1[15]&r2[2]&act_func_2_1|r1[15]&r2[3]&act_func|r1[15]&r2[3]&act_func_2_1|r1[15]&r2[4]&act_func|r1[15]&r2[4]&act_func_2_1|r1[15]&r2[5]&act_func|r1[15]&r2[5]&act_func_2_1|r1[15]&r2[6]&act_func|r1[15]&r2[6]&act_func_2_1|r1[15]&r2[7]&act_func|r1[15]&r2[7]&act_func_2_1|r1[15]&r2[8]&act_func|r1[15]&r2[8]&act_func_2_1|r1[15]&r2[9]&act_func|r1[15]&r2[9]&act_func_2_1|r1[15]&r2[10]&act_func|r1[15]&r2[10]&act_func_2_1|r1[15]&r2[11]&act_func|r1[15]&r2[11]&act_func_2_1|r1[15]&r2[12]&act_func|r1[15]&r2[12]&act_func_2_1|r1[15]&r2[13]&act_func|r1[15]&r2[13]&act_func_2_1|r1[15]&r2[14]&pow|r1[15]&r2[14]&act_func|r1[15]&r2[14]&act_func_2_1|r1[15]&r2[15]&sub|r1[15]&r2[15]&mul|r1[15]&r2[15]&pow|r1[15]&r2[15]&act_func|r1[15]&r2[15]&act_func_2_1};
endmodule
